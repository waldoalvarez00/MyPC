// Copyright 2025, Waldo Alvarez, https://pipflow.com
`timescale 1ns / 1ps

//=====================================================================
// 64-bit Unsigned Integer to IEEE 754 Extended Precision (80-bit) Converter
//
// Converts 64-bit unsigned integers (with separate sign) to 80-bit
// extended precision format.
//
// This module is designed for BCD conversion:
//   - BCD → Binary (64-bit unsigned) → FP80
//
// Features:
// - Handles unsigned 64-bit integers with separate sign bit
// - Proper normalization
// - Zero handling
// - Single-cycle operation
//=====================================================================

module FPU_UInt64_to_FP80(
    input wire clk,
    input wire reset,
    input wire enable,              // Start conversion

    // Input
    input wire [63:0] uint_in,      // 64-bit unsigned integer
    input wire        sign_in,      // Sign bit (0=positive, 1=negative)

    // Output
    output reg [79:0] fp_out,       // 80-bit floating-point
    output reg done                 // Conversion complete
);

    //=================================================================
    // Internal Registers
    //=================================================================

    reg        result_sign;
    reg [14:0] result_exp;
    reg [63:0] result_mant;
    reg [63:0] abs_value;
    reg [6:0]  shift_amount;
    integer    i;

    //=================================================================
    // Conversion Logic
    //=================================================================

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            fp_out <= 80'd0;
            done <= 1'b0;
        end else begin
            if (enable) begin
                // Handle zero
                if (uint_in == 64'd0) begin
                    fp_out <= 80'd0;  // +0.0
                    done <= 1'b1;
                end else begin
                    // Get sign and value
                    result_sign = sign_in;
                    abs_value = uint_in;

                    // Find leading 1 position (normalization)
                    shift_amount = 7'd0;
                    for (i = 63; i >= 0; i = i - 1) begin
                        if (abs_value[i] && shift_amount == 7'd0) begin
                            shift_amount = 7'd63 - i[6:0];
                        end
                    end

                    // Calculate exponent: bias + (63 - shift_amount)
                    // The integer bit will be at position 63 after shift
                    result_exp = 15'd16383 + (15'd63 - {8'd0, shift_amount});

                    // Normalize mantissa: shift so MSB is at position 63 (integer bit)
                    result_mant = abs_value << shift_amount;

                    // Pack result
                    fp_out <= {result_sign, result_exp, result_mant};
                    done <= 1'b1;
                end
            end else begin
                done <= 1'b0;
            end
        end
    end

endmodule
