// ================================================================
// Unit Test for KF8259_Interrupt_Request
// Tests edge/level triggering, freeze, and clear logic
// ================================================================

`timescale 1ns/1ps

module kf8259_interrupt_request_tb;

    // DUT signals
    logic clock;
    logic reset;
    logic level_or_edge_triggered_config;
    logic freeze;
    logic [7:0] clear_interrupt_request;
    logic [7:0] interrupt_request_pin;
    logic [7:0] interrupt_request_register;

    // Instantiate DUT
    KF8259_Interrupt_Request dut (
        .clock(clock),
        .reset(reset),
        .level_or_edge_triggered_config(level_or_edge_triggered_config),
        .freeze(freeze),
        .clear_interrupt_request(clear_interrupt_request),
        .interrupt_request_pin(interrupt_request_pin),
        .interrupt_request_register(interrupt_request_register)
    );

    // Clock generation
    initial begin
        clock = 0;
        forever #10 clock = ~clock;
    end

    // Test counters
    int test_count = 0;
    int pass_count = 0;
    int fail_count = 0;

    task check_result(input string test_name, input logic condition);
        test_count++;
        if (condition) begin
            $display("[PASS] Test %0d: %s", test_count, test_name);
            pass_count++;
        end else begin
            $display("[FAIL] Test %0d: %s", test_count, test_name);
            fail_count++;
        end
    endtask

    // Test sequence
    initial begin
        $display("================================================================");
        $display("KF8259_Interrupt_Request Unit Test");
        $display("================================================================");

        // Initialize
        reset = 1;
        level_or_edge_triggered_config = 0;  // Edge-triggered
        freeze = 0;
        clear_interrupt_request = 8'h00;
        interrupt_request_pin = 8'h00;

        repeat(5) @(posedge clock);
        reset = 0;
        repeat(2) @(posedge clock);

        // ================================================================
        // TEST 1: Edge-Triggered Mode - Rising Edge Detection
        // ================================================================
        $display("\n--- Test 1: Edge-Triggered Mode - Rising Edge ---");

        level_or_edge_triggered_config = 0;  // Edge mode
        freeze = 0;

        // Generate rising edge on IRQ0
        interrupt_request_pin[0] = 0;
        repeat(2) @(posedge clock);
        interrupt_request_pin[0] = 1;
        repeat(2) @(posedge clock);

        check_result("Edge-triggered IRQ0 latched", interrupt_request_register[0] == 1'b1);

        // Hold high - should stay latched
        repeat(5) @(posedge clock);
        check_result("Edge-triggered IRQ0 stays latched", interrupt_request_register[0] == 1'b1);

        interrupt_request_pin[0] = 0;
        repeat(2) @(posedge clock);

        // ================================================================
        // TEST 2: Edge-Triggered - Clear Request
        // ================================================================
        $display("\n--- Test 2: Edge-Triggered - Clear Request ---");

        // Trigger IRQ1
        interrupt_request_pin[1] = 0;
        repeat(2) @(posedge clock);
        interrupt_request_pin[1] = 1;
        repeat(2) @(posedge clock);

        check_result("IRQ1 latched", interrupt_request_register[1] == 1'b1);

        // Clear IRQ1
        clear_interrupt_request[1] = 1;
        @(posedge clock);
        clear_interrupt_request[1] = 0;
        @(posedge clock);

        check_result("IRQ1 cleared", interrupt_request_register[1] == 1'b0);

        interrupt_request_pin[1] = 0;
        @(posedge clock);

        // ================================================================
        // TEST 3: Edge-Triggered - Multiple Edges
        // ================================================================
        $display("\n--- Test 3: Edge-Triggered - Multiple Edges ---");

        // First edge
        interrupt_request_pin[2] = 0;
        repeat(2) @(posedge clock);
        interrupt_request_pin[2] = 1;
        repeat(2) @(posedge clock);

        check_result("First edge detected", interrupt_request_register[2] == 1'b1);

        // Clear
        clear_interrupt_request[2] = 1;
        @(posedge clock);
        clear_interrupt_request[2] = 0;
        @(posedge clock);

        // Second edge
        interrupt_request_pin[2] = 0;
        repeat(2) @(posedge clock);
        interrupt_request_pin[2] = 1;
        repeat(2) @(posedge clock);

        check_result("Second edge detected", interrupt_request_register[2] == 1'b1);

        interrupt_request_pin[2] = 0;
        clear_interrupt_request[2] = 1;
        @(posedge clock);
        clear_interrupt_request[2] = 0;
        @(posedge clock);

        // ================================================================
        // TEST 4: Level-Triggered Mode
        // ================================================================
        $display("\n--- Test 4: Level-Triggered Mode ---");

        level_or_edge_triggered_config = 1;  // Level mode
        freeze = 0;

        // Set IRQ3 high
        interrupt_request_pin[3] = 1;
        repeat(3) @(posedge clock);

        check_result("Level-triggered IRQ3 active", interrupt_request_register[3] == 1'b1);

        // Release IRQ3
        interrupt_request_pin[3] = 0;
        repeat(3) @(posedge clock);

        check_result("Level-triggered IRQ3 inactive", interrupt_request_register[3] == 1'b0);

        // ================================================================
        // TEST 5: Freeze Signal
        // ================================================================
        $display("\n--- Test 5: Freeze Signal ---");

        level_or_edge_triggered_config = 0;  // Edge mode
        freeze = 1;  // Freeze active

        // Try to trigger IRQ4 while frozen
        interrupt_request_pin[4] = 0;
        repeat(2) @(posedge clock);
        interrupt_request_pin[4] = 1;
        repeat(3) @(posedge clock);

        check_result("IRQ4 not latched while frozen", interrupt_request_register[4] == 1'b0);

        // Unfreeze
        freeze = 0;
        repeat(2) @(posedge clock);

        check_result("IRQ4 latched after unfreeze", interrupt_request_register[4] == 1'b1);

        interrupt_request_pin[4] = 0;
        clear_interrupt_request[4] = 1;
        @(posedge clock);
        clear_interrupt_request[4] = 0;
        @(posedge clock);

        // ================================================================
        // TEST 6: All IRQ Lines Simultaneously (Edge)
        // ================================================================
        $display("\n--- Test 6: All IRQ Lines Simultaneously (Edge) ---");

        level_or_edge_triggered_config = 0;
        freeze = 0;

        // Trigger all IRQs
        interrupt_request_pin = 8'h00;
        repeat(2) @(posedge clock);
        interrupt_request_pin = 8'hFF;
        repeat(3) @(posedge clock);

        check_result("All IRQs latched", interrupt_request_register == 8'hFF);

        // Clear all
        clear_interrupt_request = 8'hFF;
        @(posedge clock);
        clear_interrupt_request = 8'h00;
        @(posedge clock);

        check_result("All IRQs cleared", interrupt_request_register == 8'h00);

        interrupt_request_pin = 8'h00;
        @(posedge clock);

        // ================================================================
        // TEST 7: Selective Clear
        // ================================================================
        $display("\n--- Test 7: Selective Clear ---");

        // Trigger IRQ5, IRQ6, IRQ7
        interrupt_request_pin = 8'h00;
        repeat(2) @(posedge clock);
        interrupt_request_pin = 8'hE0;  // Bits 7, 6, 5
        repeat(3) @(posedge clock);

        check_result("IRQ5-7 latched", interrupt_request_register == 8'hE0);

        // Clear only IRQ6
        clear_interrupt_request = 8'h40;
        @(posedge clock);
        clear_interrupt_request = 8'h00;
        @(posedge clock);

        check_result("Only IRQ6 cleared", interrupt_request_register == 8'hA0);

        interrupt_request_pin = 8'h00;
        clear_interrupt_request = 8'hFF;
        @(posedge clock);
        clear_interrupt_request = 8'h00;
        @(posedge clock);

        // ================================================================
        // TEST 8: Edge Detection with Glitches
        // ================================================================
        $display("\n--- Test 8: Edge Detection with Short Pulses ---");

        level_or_edge_triggered_config = 0;
        freeze = 0;

        // Very short pulse (1 clock)
        interrupt_request_pin[0] = 0;
        @(posedge clock);
        interrupt_request_pin[0] = 1;
        @(posedge clock);
        interrupt_request_pin[0] = 0;
        repeat(2) @(posedge clock);

        check_result("Short pulse detected", interrupt_request_register[0] == 1'b1);

        clear_interrupt_request = 8'hFF;
        @(posedge clock);
        clear_interrupt_request = 8'h00;
        @(posedge clock);

        // ================================================================
        // TEST 9: Level Mode - Continuous High
        // ================================================================
        $display("\n--- Test 9: Level Mode - Continuous High ---");

        level_or_edge_triggered_config = 1;
        freeze = 0;

        // Hold IRQ1 high continuously
        interrupt_request_pin[1] = 1;
        repeat(10) @(posedge clock);

        check_result("Level mode stays active while high", interrupt_request_register[1] == 1'b1);

        interrupt_request_pin[1] = 0;
        repeat(2) @(posedge clock);

        check_result("Level mode clears when low", interrupt_request_register[1] == 1'b0);

        // ================================================================
        // TEST 10: Mode Switching
        // ================================================================
        $display("\n--- Test 10: Mode Switching (Edge to Level) ---");

        // Start in edge mode, trigger IRQ2
        level_or_edge_triggered_config = 0;
        interrupt_request_pin[2] = 0;
        repeat(2) @(posedge clock);
        interrupt_request_pin[2] = 1;
        repeat(2) @(posedge clock);

        check_result("Edge mode: IRQ2 latched", interrupt_request_register[2] == 1'b1);

        // Switch to level mode while pin still high
        level_or_edge_triggered_config = 1;
        repeat(2) @(posedge clock);

        check_result("Level mode: IRQ2 still active", interrupt_request_register[2] == 1'b1);

        // Release pin
        interrupt_request_pin[2] = 0;
        repeat(2) @(posedge clock);

        check_result("Level mode: IRQ2 cleared", interrupt_request_register[2] == 1'b0);

        // ================================================================
        // TEST 11: Reset Behavior
        // ================================================================
        $display("\n--- Test 11: Reset Behavior ---");

        // Set some IRQs
        level_or_edge_triggered_config = 0;
        interrupt_request_pin = 8'h00;
        repeat(2) @(posedge clock);
        interrupt_request_pin = 8'h55;
        repeat(3) @(posedge clock);

        // Assert reset
        reset = 1;
        repeat(2) @(posedge clock);
        reset = 0;
        repeat(2) @(posedge clock);

        check_result("Reset clears all IRQs", interrupt_request_register == 8'h00);

        interrupt_request_pin = 8'h00;
        @(posedge clock);

        // ================================================================
        // Test Summary
        // ================================================================
        $display("\n================================================================");
        $display("TEST SUMMARY");
        $display("================================================================");
        $display("Total Tests: %0d", test_count);
        $display("Passed:      %0d", pass_count);
        $display("Failed:      %0d", fail_count);
        $display("Pass Rate:   %0d%%", (pass_count * 100) / test_count);
        $display("================================================================");

        if (fail_count == 0) begin
            $display("✓✓✓ ALL TESTS PASSED ✓✓✓");
            $finish(0);
        end else begin
            $display("✗✗✗ SOME TESTS FAILED ✗✗✗");
            $finish(1);
        end
    end

    // Timeout
    initial begin
        #50000;
        $display("\n[ERROR] Testbench timeout!");
        $finish(1);
    end

endmodule
