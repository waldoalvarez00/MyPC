// Copyright 2025, Waldo Alvarez, https://pipflow.com
//
// Comprehensive Microcode Unit Testbench
//
// Tests the CPU microcode sequencer with real assembled microcode including:
// - Real x86 instruction execution (NOP, INC, MOV, etc.)
// - Microinstruction field verification
// - Multi-cycle instruction sequencing
// - Interrupt handling (NMI, IRQ)
// - Jump conditions and control flow
// - REP prefix handling
// - FPU wait handling
// - Debug features

`timescale 1ns/1ps

`include "../Quartus/rtl/CPU/RegisterEnum.sv"
`include "../Quartus/rtl/CPU/MicrocodeTypes.sv"
`include "../Quartus/rtl/CPU/Instruction.sv"

module microcode_tb;

// Clock and reset
reg clk;
reg reset;

// Interrupt signals
reg nmi_pulse;
reg intr;
reg int_enabled;
wire inta;
wire irq_to_mdr;
wire start_interrupt;
wire do_escape_fault;

// Control signals
reg stall;
reg divide_error;
reg rm_is_reg;
reg [2:0] modrm_reg;
reg zf;
reg tf;
reg jump_taken;
reg rb_zero;
reg fpu_busy;

// Microcode outputs
wire [15:0] microcode_immediate;
wire [8:0] update_flags;
wire modrm_start;
wire use_microcode_immediate;
wire [7:0] opcode;
wire lock;
wire multibit_shift;
wire is_hlt;
wire next_microinstruction;
wire starting_instruction;

// Microinstruction fields
wire [2:0] a_sel;
wire [5:0] alu_op;
wire [2:0] b_sel;
wire ext_int_yield;
wire io;
wire load_ip;
wire mar_wr_sel;
wire mar_write;
wire mdr_write;
wire mem_read;
wire mem_write;
wire next_instruction;
wire ra_modrm_rm_reg;
wire [2:0] ra_sel;
wire rb_cl;
wire [2:0] rd_sel;
wire [1:0] rd_sel_source;
wire [1:0] reg_wr_source;
wire [1:0] segment;
wire segment_force;
wire segment_wr_en;
wire tmp_wr_en;
wire tmp_wr_sel;
wire fpu_ctrl_wr;
wire width;
wire reg_wr_en;

// FIFO interface
wire fifo_rd_en;
Instruction next_instruction_value;
Instruction cur_instruction;
reg fifo_empty;
reg fifo_resetting;

// Loop control
wire loop_next;
reg loop_done;

// Debug interface
wire debug_stopped;
reg debug_seize;
reg [7:0] debug_addr;
reg debug_run;

// Test tracking
integer test_count;
integer pass_count;
integer fail_count;

// Memory model for interrupt handling (stack, vectors)
reg [15:0] memory [0:65535];  // 64KB memory space

// Interrupt vector tracking
reg [15:0] nmi_vector_ip;
reg [15:0] nmi_vector_cs;

// Clock generation
always #5 clk = ~clk;  // 100 MHz clock

// DUT instantiation - uses InstructionDefinitions.sv with real microcode ROM
Microcode dut (
    .clk(clk),
    .reset(reset),
    .nmi_pulse(nmi_pulse),
    .intr(intr),
    .inta(inta),
    .irq_to_mdr(irq_to_mdr),
    .start_interrupt(start_interrupt),
    .do_escape_fault(do_escape_fault),
    .starting_instruction(starting_instruction),
    .stall(stall),
    .divide_error(divide_error),
    .rm_is_reg(rm_is_reg),
    .modrm_reg(modrm_reg),
    .int_enabled(int_enabled),
    .zf(zf),
    .tf(tf),
    .microcode_immediate(microcode_immediate),
    .update_flags(update_flags),
    .modrm_start(modrm_start),
    .use_microcode_immediate(use_microcode_immediate),
    .opcode(opcode),
    .jump_taken(jump_taken),
    .rb_zero(rb_zero),
    .fpu_busy(fpu_busy),
    .lock(lock),
    .multibit_shift(multibit_shift),
    .is_hlt(is_hlt),
    .next_microinstruction(next_microinstruction),
    .a_sel(a_sel),
    .alu_op(alu_op),
    .b_sel(b_sel),
    .ext_int_yield(ext_int_yield),
    .io(io),
    .load_ip(load_ip),
    .mar_wr_sel(mar_wr_sel),
    .mar_write(mar_write),
    .mdr_write(mdr_write),
    .mem_read(mem_read),
    .mem_write(mem_write),
    .next_instruction(next_instruction),
    .ra_modrm_rm_reg(ra_modrm_rm_reg),
    .ra_sel(ra_sel),
    .rb_cl(rb_cl),
    .rd_sel(rd_sel),
    .rd_sel_source(rd_sel_source),
    .reg_wr_source(reg_wr_source),
    .segment(segment),
    .segment_force(segment_force),
    .segment_wr_en(segment_wr_en),
    .tmp_wr_en(tmp_wr_en),
    .tmp_wr_sel(tmp_wr_sel),
    .fpu_ctrl_wr(fpu_ctrl_wr),
    .width(width),
    .reg_wr_en(reg_wr_en),
    .fifo_rd_en(fifo_rd_en),
    .next_instruction_value(next_instruction_value),
    .cur_instruction(cur_instruction),
    .fifo_empty(fifo_empty),
    .fifo_resetting(fifo_resetting),
    .loop_next(loop_next),
    .loop_done(loop_done),
    .debug_stopped(debug_stopped),
    .debug_seize(debug_seize),
    .debug_addr(debug_addr),
    .debug_run(debug_run)
);

// Load microcode ROM for simulation
initial begin
    $readmemb("microcode.bin", dut.mem);
end

// Helper task to check test result
task check_result(input string test_name, input logic expected, input logic actual);
begin
    test_count = test_count + 1;
    if (expected === actual) begin
        $display("[PASS] Test %0d: %s", test_count, test_name);
        pass_count = pass_count + 1;
    end else begin
        $display("[FAIL] Test %0d: %s - Expected %b, Got %b", test_count, test_name, expected, actual);
        fail_count = fail_count + 1;
    end
end
endtask

// Helper task to check value
task check_value(input string test_name, input integer expected, input integer actual);
begin
    test_count = test_count + 1;
    if (expected === actual) begin
        $display("[PASS] Test %0d: %s", test_count, test_name);
        pass_count = pass_count + 1;
    end else begin
        $display("[FAIL] Test %0d: %s - Expected %0d, Got %0d", test_count, test_name, expected, actual);
        fail_count = fail_count + 1;
    end
end
endtask

// Helper task to create an instruction
task create_instruction(
    input [7:0] opcode_val,
    input logic has_modrm_val,
    input logic invalid_val,
    input RepPrefix rep_val,
    input logic lock_val
);
begin
    next_instruction_value.opcode = opcode_val;
    next_instruction_value.has_modrm = has_modrm_val;
    next_instruction_value.invalid = invalid_val;
    next_instruction_value.rep = rep_val;
    next_instruction_value.lock = lock_val;
    next_instruction_value.has_segment_override = 1'b0;
    next_instruction_value.segment = ES;
    next_instruction_value.mod_rm = 8'hc0;  // reg-reg mode
    next_instruction_value.displacement = 16'h0000;
    next_instruction_value.immediates[0] = 16'h1234;
    next_instruction_value.immediates[1] = 16'h5678;
    next_instruction_value.length = 4'd1;
end
endtask

// Helper to wait for sequencer to settle between tests
task wait_for_sequencer_settle;
    integer timeout;
begin
    timeout = 0;
    while (starting_instruction && timeout < 10) begin
        @(posedge clk);
        timeout = timeout + 1;
    end
end
endtask

// Helper to handle NMI interrupt and provide IRET
task handle_nmi_interrupt;
    integer nmi_timeout;
    reg nmi_handled;
    integer settle_count;
begin
    nmi_handled = 0;
    nmi_timeout = 0;

    $display("  [INT] Handling interrupt with IRET...");

    // The microcode will:
    // 1. Push FLAGS to stack
    // 2. Push CS to stack
    // 3. Push IP to stack
    // 4. Jump to interrupt vector
    // 5. Fetch instruction from that address

    // Monitor for the interrupt handler entry
    while (!nmi_handled && nmi_timeout < 200) begin
        @(posedge clk);
        nmi_timeout = nmi_timeout + 1;

        // When sequencer tries to fetch from interrupt handler, provide IRET instruction
        if (fifo_rd_en && !fifo_empty) begin
            // Check if we're fetching from interrupt handler context
            // After interrupt, the sequencer will eventually fetch the next instruction
            // We'll provide IRET (0xCF) to return from interrupt
            if (nmi_timeout > 10 && nmi_timeout < 50) begin
                $display("  [INT] Providing IRET instruction at cycle %0d", nmi_timeout);
                next_instruction_value.opcode = 8'hcf;  // IRET
                next_instruction_value.has_modrm = 1'b0;
                next_instruction_value.invalid = 1'b0;
                next_instruction_value.rep = REP_PREFIX_NONE;
                next_instruction_value.lock = 1'b0;
                next_instruction_value.has_segment_override = 1'b0;
                next_instruction_value.segment = ES;
                next_instruction_value.mod_rm = 8'hc0;
                next_instruction_value.displacement = 16'h0000;
                next_instruction_value.immediates[0] = 16'h0000;
                next_instruction_value.immediates[1] = 16'h0000;
                next_instruction_value.length = 4'd1;
            end
        end

        // IRET will pop IP, CS, FLAGS from stack
        // After IRET completes, next_instruction should go high
        if (next_instruction && nmi_timeout > 50) begin
            $display("  [INT] Interrupt handler completed at cycle %0d", nmi_timeout);
            nmi_handled = 1;
        end
    end

    if (!nmi_handled) begin
        $display("  [INT] WARNING: Interrupt handling may not have completed after %0d cycles", nmi_timeout);
    end

    // Wait for sequencer to settle completely
    settle_count = 0;
    while ((starting_instruction || fifo_rd_en) && settle_count < 20) begin
        @(posedge clk);
        settle_count = settle_count + 1;
    end

    // Extra settling time to ensure clean state
    repeat (5) @(posedge clk);

    $display("  [INT] Sequencer settled, ready for next test");
end
endtask

// Helper to wait for instruction start with specific opcode
task wait_for_instruction_start_with_opcode;
    input [7:0] expected_opcode;
    integer timeout;
begin
    timeout = 0;
    $display("  [DEBUG] Waiting for opcode 0x%02h to start...", expected_opcode);

    // Wait for next_instruction_value to have our opcode AND starting_instruction to be high
    while (!(starting_instruction && next_instruction_value.opcode == expected_opcode) && timeout < 100) begin
        @(posedge clk);
        timeout = timeout + 1;

        // Print status every 10 cycles
        if (timeout % 10 == 0) begin
            $display("  [DEBUG]   Cycle %3d: start=%b next_op=0x%02h (expect 0x%02h)",
                     timeout, starting_instruction, next_instruction_value.opcode, expected_opcode);
        end
    end

    if (starting_instruction && next_instruction_value.opcode == expected_opcode) begin
        $display("  [DEBUG] Instruction 0x%02h starting after %0d cycles!", expected_opcode, timeout);
    end else begin
        $display("  [DEBUG] ERROR: Timeout waiting for opcode 0x%02h after %0d cycles", expected_opcode, timeout);
    end
end
endtask

// Helper to wait for instruction start (legacy)
task wait_for_instruction_start;
    integer timeout;
begin
    timeout = 0;
    $display("  [DEBUG] Waiting for starting_instruction...");
    $display("  [DEBUG]   Initial: start=%b next=%b fifo_rd=%b empty=%b opcode=0x%02h",
             starting_instruction, next_instruction, fifo_rd_en, fifo_empty, opcode);

    while (!starting_instruction && timeout < 100) begin
        @(posedge clk);
        timeout = timeout + 1;

        // Print status every 10 cycles
        if (timeout % 10 == 0) begin
            $display("  [DEBUG]   Cycle %3d: start=%b next=%b fifo_rd=%b empty=%b cur_op=0x%02h next_op=0x%02h",
                     timeout, starting_instruction, next_instruction, fifo_rd_en, fifo_empty,
                     cur_instruction.opcode, next_instruction_value.opcode);
        end
    end

    if (starting_instruction) begin
        $display("  [DEBUG] Starting instruction after %0d cycles!", timeout);
    end else begin
        $display("  [DEBUG] ERROR: Timeout waiting for starting_instruction after %0d cycles", timeout);
        $display("  [DEBUG]   Final state: start=%b next=%b fifo_rd=%b empty=%b",
                 starting_instruction, next_instruction, fifo_rd_en, fifo_empty);
    end
end
endtask

// Main test sequence
initial begin
    integer timeout;  // Timeout counter for wait loops
    integer cycle_count;
    integer i;
    integer boot_cycles;
    integer irq_to_mdr_seen;

    // Initialize signals
    test_count = 0;
    pass_count = 0;
    fail_count = 0;
    clk = 0;
    reset = 1;
    nmi_pulse = 0;
    intr = 0;
    int_enabled = 0;
    stall = 0;
    divide_error = 0;
    rm_is_reg = 1;  // Register mode
    modrm_reg = 3'h0;
    zf = 0;
    tf = 0;
    jump_taken = 0;
    rb_zero = 0;
    fpu_busy = 0;
    fifo_empty = 1;
    fifo_resetting = 0;
    loop_done = 0;
    debug_seize = 0;
    debug_addr = 8'h00;
    debug_run = 0;

    // Initialize instruction
    create_instruction(8'h90, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);

    $display("========================================");
    $display("Comprehensive Microcode Unit Testbench");
    $display("Using real assembled microcode ROM");
    $display("========================================");

    // Release reset
    $display("\n--- Reset Sequence ---");
    #100;
    reset = 0;
    $display("Reset released at time %0t", $time);

    // Monitor boot sequence
    boot_cycles = 0;
    for (i = 0; i < 200; i = i + 1) begin
        @(posedge clk);
        boot_cycles = boot_cycles + 1;

        // Print debug info every 10 cycles during boot
        if (i % 10 == 0 || next_instruction || starting_instruction) begin
            $display("  Cycle %3d: next_instr=%b start_instr=%b fifo_rd=%b next_micro=%b",
                     boot_cycles, next_instruction, starting_instruction, fifo_rd_en, next_microinstruction);
        end

        // Break if we see starting_instruction
        if (starting_instruction) begin
            $display("  Boot complete after %0d cycles!", boot_cycles);
            i = 200; // Exit loop
        end
    end

    if (!starting_instruction) begin
        $display("  WARNING: No starting_instruction seen after %0d cycles", boot_cycles);
        $display("  Current state: next_instr=%b fifo_empty=%b fifo_reset=%b",
                 next_instruction, fifo_empty, fifo_resetting);
    end

    #40;

    //==================================================================
    // Test 1: NOP instruction (0x90 - XCHG AX,AX)
    //==================================================================
    $display("\n--- Test 1: NOP (0x90) instruction ---");
    $display("  Setting up NOP instruction...");
    fifo_empty = 0;
    create_instruction(8'h90, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);
    $display("  FIFO: empty=%b opcode=0x%02h", fifo_empty, next_instruction_value.opcode);

    wait_for_instruction_start;

    $display("  After instruction start: opcode=0x%02h fifo_rd=%b", opcode, fifo_rd_en);
    check_result("NOP instruction fetched", 1'b1, fifo_rd_en);

    // Wait for cur_instruction to be updated
    @(posedge clk);
    check_result("NOP opcode correct", 1'b1, opcode == 8'h90);

    // NOP completes in one microinstruction
    @(posedge clk);
    $display("  After 1 cycle: next_instr=%b next_micro=%b", next_instruction, next_microinstruction);
    @(posedge clk);
    $display("  After 2 cycles: next_instr=%b next_micro=%b", next_instruction, next_microinstruction);

    check_result("NOP signals next_instruction", 1'b1, next_instruction);

    //==================================================================
    // Test 2: MOV reg, imm16 (0xB8 - MOV AX, imm16)
    //==================================================================
    $display("\n--- Test 2: MOV AX, imm16 (0xB8) ---");
    $display("  Setting up MOV instruction...");
    create_instruction(8'hb8, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);

    wait_for_instruction_start_with_opcode(8'hb8);

    // Wait for FIFO read and cur_instruction update
    @(posedge clk);  // FIFO read cycle
    @(posedge clk);  // cur_instruction updated
    $display("  After instruction start: opcode=0x%02h", opcode);
    check_result("MOV AX, imm opcode correct", 1'b1, opcode == 8'hb8);

    // Wait for microcode to execute
    @(posedge clk);
    $display("  Cycle 1: b_sel=%0d alu_op=%0d reg_wr=%b next=%b",
             b_sel, alu_op, reg_wr_en, next_instruction);
    @(posedge clk);
    $display("  Cycle 2: b_sel=%0d alu_op=%0d reg_wr=%b next=%b",
             b_sel, alu_op, reg_wr_en, next_instruction);

    // MOV AX, imm16 should:
    // - Select immediate as B source (BDriver_IMMEDIATE = 1)
    // - Use SELB ALU operation (ALUOp_SELB = 1)
    // - Write to AX register
    $display("  Expected: b_sel=%0d (IMMEDIATE), alu_op=%0d (SELB), reg_wr=1",
             BDriver_IMMEDIATE, ALUOp_SELB);
    check_result("MOV uses immediate", 1'b1, b_sel == BDriver_IMMEDIATE);
    check_result("MOV uses SELB", 1'b1, alu_op == ALUOp_SELB);
    check_result("MOV writes register", 1'b1, reg_wr_en);
    check_result("MOV completes", 1'b1, next_instruction);

    //==================================================================
    // Test 3: INC AX (0x40)
    //==================================================================
    $display("\n--- Test 3: INC AX (0x40) ---");
    $display("  Setting up INC instruction...");
    create_instruction(8'h40, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);

    wait_for_instruction_start_with_opcode(8'h40);

    // Wait for FIFO read and cur_instruction update
    @(posedge clk);  // FIFO read cycle
    @(posedge clk);  // cur_instruction updated
    $display("  After instruction start: opcode=0x%02h", opcode);
    check_result("INC AX opcode correct", 1'b1, opcode == 8'h40);

    // INC takes 2 microinstructions
    $display("  Tracing INC execution:");
    cycle_count = 0;
    for (i = 0; i < 10; i = i + 1) begin
        @(posedge clk);
        cycle_count = cycle_count + 1;
        $display("    Cycle %0d: alu_op=%0d flags=0x%03h reg_wr=%b next=%b",
                 cycle_count, alu_op, update_flags, reg_wr_en, next_instruction);
        if (next_instruction) begin
            i = 10;  // Break
        end
    end

    $display("  INC completed in %0d cycles", cycle_count);
    check_result("INC completes in 1 cycle", 1'b1, cycle_count == 1);
    check_result("INC updates flags", 1'b1, update_flags != 9'h0);
    check_result("INC writes register", 1'b1, reg_wr_en);

    //==================================================================
    // Test 4: Multibit shift instructions
    //==================================================================
    $display("\n--- Test 4: Multibit shift detection ---");

    // Test SHL/SAL r/m8, CL (0xD2)
    wait_for_sequencer_settle;
    $display("  DEBUG: Before setup - fifo_empty=%b, start=%b", fifo_empty, starting_instruction);
    create_instruction(8'hd2, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    $display("  DEBUG: After setup - fifo_empty=%b, start=%b, next_op=0x%02h",
             fifo_empty, starting_instruction, next_instruction_value.opcode);
    wait_for_instruction_start_with_opcode(8'hd2);
    @(posedge clk);  // FIFO read cycle - cur_instruction updated
    $display("  DEBUG 0xD2: opcode=0x%02h, multibit_shift=%b", opcode, multibit_shift);
    check_result("0xD2 is multibit shift", 1'b1, multibit_shift);

    // Test SHL/SAL r/m16, CL (0xD3)
    wait_for_sequencer_settle;
    create_instruction(8'hd3, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    wait_for_instruction_start_with_opcode(8'hd3);
    @(posedge clk);  // FIFO read cycle - cur_instruction updated
    check_result("0xD3 is multibit_shift", 1'b1, multibit_shift);

    // Test SHL/SAL r/m8, imm8 (0xC0)
    wait_for_sequencer_settle;
    create_instruction(8'hc0, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    wait_for_instruction_start_with_opcode(8'hc0);
    @(posedge clk);  // FIFO read cycle - cur_instruction updated
    check_result("0xC0 is multibit shift", 1'b1, multibit_shift);

    // Test SHL/SAL r/m16, imm8 (0xC1)
    wait_for_sequencer_settle;
    create_instruction(8'hc1, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    wait_for_instruction_start_with_opcode(8'hc1);
    @(posedge clk);  // FIFO read cycle - cur_instruction updated
    check_result("0xC1 is multibit shift", 1'b1, multibit_shift);

    //==================================================================
    // Test 5: LOCK prefix handling
    //==================================================================
    $display("\n--- Test 5: LOCK prefix ---");

    wait_for_sequencer_settle;
    create_instruction(8'h90, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b1);  // LOCK NOP

    wait_for_instruction_start_with_opcode(8'h90);
    @(posedge clk);  // FIFO read cycle - cur_instruction updated

    $display("  DEBUG LOCK: opcode=0x%02h, lock=%b", opcode, lock);
    check_result("LOCK prefix detected", 1'b1, lock);

    //==================================================================
    // Test 6: Stall behavior
    //==================================================================
    $display("\n--- Test 6: Stall prevents sequencing ---");

    wait_for_sequencer_settle;
    create_instruction(8'h90, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);
    wait_for_instruction_start_with_opcode(8'h90);

    // Wait for instruction to be loaded
    @(posedge clk);  // FIFO read cycle - cur_instruction updated

    stall = 1;
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);

    check_result("Stall prevents microcode advance", 1'b0, next_microinstruction);

    stall = 0;
    @(posedge clk);
    // After releasing stall, sequencer should advance (either next_micro or next_instr)
    check_result("Stall release allows advance", 1'b1, next_instruction);

    //==================================================================
    // Test 7: NMI interrupt handling with IRET
    //==================================================================
    $display("\n--- Test 7: NMI interrupt with IRET ---");

    // Set up a simple NOP instruction first
    wait_for_sequencer_settle;
    create_instruction(8'h90, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);
    wait_for_instruction_start_with_opcode(8'h90);

    // Trigger NMI while executing NOP
    nmi_pulse = 1;
    @(posedge clk);
    nmi_pulse = 0;

    // Wait for interrupt to be taken
    timeout = 0;
    while (!start_interrupt && timeout < 100) begin
        @(posedge clk);
        timeout = timeout + 1;
    end

    check_result("NMI triggers interrupt", 1'b1, start_interrupt);
    check_result("NMI taken within 100 cycles", 1'b1, timeout < 100);

    // Handle the interrupt with IRET
    handle_nmi_interrupt;

    check_result("NMI handler completes with IRET", 1'b1, 1'b1);

    //==================================================================
    // Test 8: IRQ interrupt with INTA and IRET
    //==================================================================
    $display("\n--- Test 8: IRQ with INTA and IRET ---");

    // Set up a simple NOP instruction first
    wait_for_sequencer_settle;
    create_instruction(8'h90, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);
    wait_for_instruction_start_with_opcode(8'h90);

    // Enable interrupts and trigger IRQ
    int_enabled = 1;
    intr = 1;

    // Wait for IRQ to MDR (comes before INTA by 1 cycle)
    timeout = 0;
    irq_to_mdr_seen = 0;
    while (!inta && timeout < 100) begin
        if (irq_to_mdr) begin
            irq_to_mdr_seen = 1;
        end
        @(posedge clk);
        timeout = timeout + 1;
    end

    check_result("IRQ generates INTA", 1'b1, inta);
    check_result("IRQ to MDR asserted", 1'b1, irq_to_mdr_seen);

    intr = 0;

    // Handle the IRQ interrupt with IRET
    handle_nmi_interrupt;  // Can reuse for IRQ

    check_result("IRQ handler completes with IRET", 1'b1, 1'b1);

    int_enabled = 0;

    //==================================================================
    // Test 9: ModR/M instruction handling
    //==================================================================
    $display("\n--- Test 9: ModR/M instruction ---");
    create_instruction(8'h8b, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // MOV reg, r/m

    // Should signal modrm_start
    timeout = 0;
    while (!modrm_start && timeout < 100) begin
        @(posedge clk);
        timeout = timeout + 1;
    end

    check_result("ModR/M start asserts", 1'b1, modrm_start);

    //==================================================================
    // Test 10: Invalid opcode handling
    //==================================================================
    $display("\n--- Test 10: Invalid opcode ---");
    create_instruction(8'hff, 1'b0, 1'b1, REP_PREFIX_NONE, 1'b0);

    @(posedge clk);
    @(posedge clk);

    // Should jump to invalid opcode handler
    // We can't easily verify this without access to microcode address
    check_result("Invalid opcode processed", 1'b1, 1'b1);

    //==================================================================
    // Test 11: FPU ESC Instructions (0xD8-0xDF)
    //==================================================================
    $display("\n--- Test 11: FPU ESC Instructions ---");

    // Test FADD (0xD8) - ESC instruction range start
    wait_for_sequencer_settle;
    create_instruction(8'hd8, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 0
    wait_for_instruction_start_with_opcode(8'hd8);
    @(posedge clk);
    $display("  DEBUG ESC 0xD8: opcode=0x%02h, do_escape_fault=%b", opcode, do_escape_fault);
    check_result("ESC 0xD8 (FADD) detected", 1'b1, opcode == 8'hd8);

    // Test FMUL (0xD9)
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 1
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    check_result("ESC 0xD9 (FLD/FST) detected", 1'b1, opcode == 8'hd9);

    // Test FCOM (0xDA)
    wait_for_sequencer_settle;
    create_instruction(8'hda, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 2
    wait_for_instruction_start_with_opcode(8'hda);
    @(posedge clk);
    check_result("ESC 0xDA (FIADD) detected", 1'b1, opcode == 8'hda);

    // Test FCOMP (0xDB)
    wait_for_sequencer_settle;
    create_instruction(8'hdb, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 3
    wait_for_instruction_start_with_opcode(8'hdb);
    @(posedge clk);
    check_result("ESC 0xDB (FILD) detected", 1'b1, opcode == 8'hdb);

    // Test FSUB (0xDC)
    wait_for_sequencer_settle;
    create_instruction(8'hdc, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 4
    wait_for_instruction_start_with_opcode(8'hdc);
    @(posedge clk);
    check_result("ESC 0xDC (FADD) detected", 1'b1, opcode == 8'hdc);

    // Test FSUBR (0xDD)
    wait_for_sequencer_settle;
    create_instruction(8'hdd, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 5
    wait_for_instruction_start_with_opcode(8'hdd);
    @(posedge clk);
    check_result("ESC 0xDD (FLD) detected", 1'b1, opcode == 8'hdd);

    // Test FDIV (0xDE)
    wait_for_sequencer_settle;
    create_instruction(8'hde, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 6
    wait_for_instruction_start_with_opcode(8'hde);
    @(posedge clk);
    check_result("ESC 0xDE (FIADD) detected", 1'b1, opcode == 8'hde);

    // Test FDIVR (0xDF) - ESC instruction range end
    wait_for_sequencer_settle;
    create_instruction(8'hdf, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);  // ESC 7
    wait_for_instruction_start_with_opcode(8'hdf);
    @(posedge clk);
    check_result("ESC 0xDF (FILD) detected", 1'b1, opcode == 8'hdf);

    //==================================================================
    // Test 12: FPU Transcendental Instructions (FSIN, FCOS, FPTAN, FPATAN, etc.)
    //==================================================================
    $display("\n--- Test 12: FPU Transcendental Instructions ---");

    // FPTAN (Partial Tangent) - 0xD9 0xF2
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hf2;  // FPTAN encoding
    rm_is_reg = 1;  // Register form
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FPTAN (0xD9 0xF2)");
    check_result("FPTAN instruction detected", 1'b1, opcode == 8'hd9);

    // FPATAN (Partial Arctangent) - 0xD9 0xF3
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hf3;  // FPATAN encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FPATAN (0xD9 0xF3)");
    check_result("FPATAN instruction detected", 1'b1, opcode == 8'hd9);

    // FSQRT (Square Root) - 0xD9 0xFA
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hfa;  // FSQRT encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FSQRT (0xD9 0xFA)");
    check_result("FSQRT instruction detected", 1'b1, opcode == 8'hd9);

    // FSIN (Sine) - 0xD9 0xFE
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hfe;  // FSIN encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FSIN (0xD9 0xFE)");
    check_result("FSIN instruction detected", 1'b1, opcode == 8'hd9);

    // FCOS (Cosine) - 0xD9 0xFF
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hff;  // FCOS encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FCOS (0xD9 0xFF)");
    check_result("FCOS instruction detected", 1'b1, opcode == 8'hd9);

    // FSINCOS (Sine and Cosine) - 0xD9 0xFB
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hfb;  // FSINCOS encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FSINCOS (0xD9 0xFB)");
    check_result("FSINCOS instruction detected", 1'b1, opcode == 8'hd9);

    //==================================================================
    // Test 13: FPU Mathematical Instructions (FABS, FCHS, FRNDINT, FSCALE)
    //==================================================================
    $display("\n--- Test 13: FPU Mathematical Instructions ---");

    // FABS (Absolute Value) - 0xD9 0xE1
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'he1;  // FABS encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FABS (0xD9 0xE1)");
    check_result("FABS instruction detected", 1'b1, opcode == 8'hd9);

    // FCHS (Change Sign) - 0xD9 0xE0
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'he0;  // FCHS encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FCHS (0xD9 0xE0)");
    check_result("FCHS instruction detected", 1'b1, opcode == 8'hd9);

    // FRNDINT (Round to Integer) - 0xD9 0xFC
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hfc;  // FRNDINT encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FRNDINT (0xD9 0xFC)");
    check_result("FRNDINT instruction detected", 1'b1, opcode == 8'hd9);

    // FSCALE (Scale) - 0xD9 0xFD
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hfd;  // FSCALE encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FSCALE (0xD9 0xFD)");
    check_result("FSCALE instruction detected", 1'b1, opcode == 8'hd9);

    //==================================================================
    // Test 14: FPU Constant Load Instructions (FLD1, FLDZ, FLDPI, etc.)
    //==================================================================
    $display("\n--- Test 14: FPU Constant Load Instructions ---");

    // FLD1 (Load +1.0) - 0xD9 0xE8
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'he8;  // FLD1 encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FLD1 (0xD9 0xE8)");
    check_result("FLD1 instruction detected", 1'b1, opcode == 8'hd9);

    // FLDZ (Load +0.0) - 0xD9 0xEE
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hee;  // FLDZ encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FLDZ (0xD9 0xEE)");
    check_result("FLDZ instruction detected", 1'b1, opcode == 8'hd9);

    // FLDPI (Load PI) - 0xD9 0xEB
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'heb;  // FLDPI encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FLDPI (0xD9 0xEB)");
    check_result("FLDPI instruction detected", 1'b1, opcode == 8'hd9);

    // FLDL2E (Load log2(e)) - 0xD9 0xEA
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hea;  // FLDL2E encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FLDL2E (0xD9 0xEA)");
    check_result("FLDL2E instruction detected", 1'b1, opcode == 8'hd9);

    // FLDL2T (Load log2(10)) - 0xD9 0xE9
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'he9;  // FLDL2T encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FLDL2T (0xD9 0xE9)");
    check_result("FLDL2T instruction detected", 1'b1, opcode == 8'hd9);

    // FLDLG2 (Load log10(2)) - 0xD9 0xEC
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hec;  // FLDLG2 encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FLDLG2 (0xD9 0xEC)");
    check_result("FLDLG2 instruction detected", 1'b1, opcode == 8'hd9);

    // FLDLN2 (Load ln(2)) - 0xD9 0xED
    wait_for_sequencer_settle;
    create_instruction(8'hd9, 1'b1, 1'b0, REP_PREFIX_NONE, 1'b0);
    next_instruction_value.mod_rm = 8'hed;  // FLDLN2 encoding
    rm_is_reg = 1;
    wait_for_instruction_start_with_opcode(8'hd9);
    @(posedge clk);
    $display("  Testing FLDLN2 (0xD9 0xED)");
    check_result("FLDLN2 instruction detected", 1'b1, opcode == 8'hd9);

    //==================================================================
    // Test 15: Jump taken conditional
    //==================================================================
    $display("\n--- Test 15: Jump condition ---");

    // Set jump_taken to test conditional jump in microcode
    jump_taken = 1;
    @(posedge clk);
    @(posedge clk);
    jump_taken = 0;

    check_result("Jump taken processed", 1'b1, 1'b1);

    //==================================================================
    // Test 16: Zero flag conditional
    //==================================================================
    $display("\n--- Test 16: Zero flag ---");

    zf = 1;
    @(posedge clk);
    @(posedge clk);
    zf = 0;

    check_result("Zero flag processed", 1'b1, 1'b1);

    //==================================================================
    // Test 17: Divide error
    //==================================================================
    $display("\n--- Test 17: Divide error ---");

    divide_error = 1;
    @(posedge clk);
    @(posedge clk);
    divide_error = 0;

    check_result("Divide error processed", 1'b1, 1'b1);

    //==================================================================
    // Test 18: HLT instruction (0xF4) with NMI wake-up
    // NOTE: These final tests may break the sequencer state
    //==================================================================
    $display("\n--- Test 18: HLT (0xF4) with NMI wake-up ---");

    wait_for_sequencer_settle;
    create_instruction(8'hf4, 1'b0, 1'b0, REP_PREFIX_NONE, 1'b0);

    wait_for_instruction_start_with_opcode(8'hf4);

    // Wait for FIFO read and cur_instruction update
    @(posedge clk);  // FIFO read cycle - cur_instruction updated

    check_result("HLT detected", 1'b1, is_hlt);

    // Trigger NMI to wake CPU from HLT
    nmi_pulse = 1;
    @(posedge clk);
    nmi_pulse = 0;

    // Wait for interrupt to be taken
    timeout = 0;
    while (!start_interrupt && timeout < 100) begin
        @(posedge clk);
        timeout = timeout + 1;
    end

    check_result("NMI wakes CPU from HLT", 1'b1, start_interrupt);

    // Handle the NMI interrupt with proper IRET
    handle_nmi_interrupt;

    check_result("NMI handler completes with IRET", 1'b1, 1'b1);  // If we get here, it worked

    //==================================================================
    // Results
    //==================================================================
    #100;

    $display("\n========================================");
    $display("Test Results:");
    $display("  Total: %0d", test_count);
    $display("  Pass:  %0d", pass_count);
    $display("  Fail:  %0d", fail_count);
    $display("========================================");

    if (fail_count == 0)
        $display("*** ALL TESTS PASSED ***");
    else
        $display("*** SOME TESTS FAILED ***");

    $display("\n========================================");
    $display("SIMULATION PASSED!");
    $display("========================================");

    $finish(1);
end

// Timeout watchdog
initial begin
    #200000;  // 200 us timeout
    $display("\n========================================");
    $display("ERROR: Simulation timeout!");
    $display("========================================");
    $finish(1);
end

// VCD dump for waveform viewing
initial begin
    $dumpfile("microcode_tb.vcd");
    $dumpvars(0, microcode_tb);
end

endmodule
