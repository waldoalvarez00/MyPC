// Copyright 2025, Waldo Alvarez, https://pipflow.com
`timescale 1ns / 1ps

//=====================================================================
// Unified Format Converter for 8087 FPU
//
// Consolidates 12+ format conversion modules into a single parameterized
// unit with mode selection.
//
// Supported Conversions:
//   - FP32 ↔ FP80
//   - FP64 ↔ FP80
//   - Int16 ↔ FP80
//   - Int32 ↔ FP80
//   - UInt64 ↔ FP80
//
// Benefits:
//   - ~60% area reduction vs. separate modules
//   - Shared rounding, normalization, and special value logic
//   - Single-cycle operation for all modes
//
// Area Savings: ~1000 lines (12 modules × 133 avg → 600 lines unified)
//=====================================================================

module FPU_Format_Converter_Unified(
    input wire clk,
    input wire reset,
    input wire enable,              // Start conversion

    // Mode selection (4 bits = 16 modes)
    input wire [3:0] mode,          // See MODE_* parameters below

    // Input ports (only relevant port is used per mode)
    input wire [79:0] fp80_in,      // FP80 input
    input wire [63:0] fp64_in,      // FP64 input
    input wire [31:0] fp32_in,      // FP32 input
    input wire [63:0] uint64_in,    // UInt64 input
    input wire [31:0] int32_in,     // Int32 input (sign-extended)
    input wire [15:0] int16_in,     // Int16 input (sign-extended)
    input wire [63:0] fixed64_in,   // Q2.62 fixed-point input (signed)
    input wire        uint64_sign,  // Sign for UInt64→FP80 (BCD)

    // Rounding mode (for FP80→narrower conversions)
    input wire [1:0] rounding_mode, // 00=nearest, 01=down, 10=up, 11=truncate

    // Output ports (only relevant port is valid per mode)
    output reg [79:0] fp80_out,     // FP80 output
    output reg [63:0] fp64_out,     // FP64 output
    output reg [31:0] fp32_out,     // FP32 output
    output reg [63:0] uint64_out,   // UInt64 output
    output reg [31:0] int32_out,    // Int32 output
    output reg [15:0] int16_out,    // Int16 output
    output reg [63:0] fixed64_out,  // Q2.62 fixed-point output (signed)
    output reg        uint64_sign_out, // Sign output for FP80→UInt64 (BCD)

    // Status
    output reg done,                // Conversion complete

    // Exception flags
    output reg flag_invalid,        // Invalid operation (NaN)
    output reg flag_overflow,       // Result overflow
    output reg flag_underflow,      // Result underflow
    output reg flag_inexact         // Result not exact (rounded)
);

    //=================================================================
    // Mode Definitions
    //=================================================================

    localparam MODE_FP32_TO_FP80  = 4'd0;
    localparam MODE_FP64_TO_FP80  = 4'd1;
    localparam MODE_FP80_TO_FP32  = 4'd2;
    localparam MODE_FP80_TO_FP64  = 4'd3;
    localparam MODE_INT16_TO_FP80 = 4'd4;
    localparam MODE_INT32_TO_FP80 = 4'd5;
    localparam MODE_FP80_TO_INT16 = 4'd6;
    localparam MODE_FP80_TO_INT32 = 4'd7;
    localparam MODE_UINT64_TO_FP80 = 4'd8;
    localparam MODE_FP80_TO_UINT64 = 4'd9;
    localparam MODE_FP80_TO_FIXED64 = 4'd10;  // FP80 → Q2.62 fixed-point for CORDIC
    localparam MODE_FIXED64_TO_FP80 = 4'd11;  // Q2.62 fixed-point → FP80 for CORDIC
    // Modes 12-15 reserved for future use (BCD, FP16, etc.)

    //=================================================================
    // Unpacked Components (shared across all formats)
    //=================================================================

    reg        src_sign;
    reg [14:0] src_exp;
    reg [63:0] src_mant;
    reg signed [16:0] src_exp_unbiased;

    reg        dst_sign;
    reg [14:0] dst_exp;
    reg [63:0] dst_mant;

    //=================================================================
    // Working Registers
    //=================================================================

    reg [6:0]  shift_amount;
    reg [63:0] shifted_mant;
    reg [63:0] abs_int_value;
    reg signed [63:0] signed_int_value;
    reg        round_up;
    reg        is_special;
    reg        is_zero;
    reg        is_inf;
    reg        is_nan;

    integer i;

    //=================================================================
    // Main Conversion Logic
    //=================================================================

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            fp80_out <= 80'd0;
            fp64_out <= 64'd0;
            fp32_out <= 32'd0;
            uint64_out <= 64'd0;
            int32_out <= 32'd0;
            int16_out <= 16'd0;
            fixed64_out <= 64'd0;
            uint64_sign_out <= 1'b0;
            done <= 1'b0;
            flag_invalid <= 1'b0;
            flag_overflow <= 1'b0;
            flag_underflow <= 1'b0;
            flag_inexact <= 1'b0;
        end else begin
            if (enable) begin
                // Clear flags
                flag_invalid = 1'b0;
                flag_overflow = 1'b0;
                flag_underflow = 1'b0;
                flag_inexact = 1'b0;

                case (mode)
                    //=============================================
                    // FP32 → FP80
                    //=============================================
                    MODE_FP32_TO_FP80: begin
                        // Unpack FP32
                        src_sign = fp32_in[31];
                        src_exp = {7'd0, fp32_in[30:23]};
                        src_mant = {fp32_in[22:0], 41'd0};  // Fraction only

                        dst_sign = src_sign;

                        // Handle special values
                        if (fp32_in[30:23] == 8'd0) begin
                            // Zero or denormalized
                            if (fp32_in[22:0] == 23'd0) begin
                                // ±0
                                dst_exp = 15'd0;
                                dst_mant = 64'd0;
                            end else begin
                                // Denormalized: normalize for FP80
                                shift_amount = 7'd0;
                                for (i = 22; i >= 0; i = i - 1) begin
                                    if (fp32_in[i] && shift_amount == 7'd0)
                                        shift_amount = 7'd22 - i[6:0];
                                end
                                dst_exp = 15'd16383 - 15'd126 - {8'd0, shift_amount};
                                dst_mant = src_mant << (shift_amount + 7'd1);
                            end
                        end else if (fp32_in[30:23] == 8'd255) begin
                            // ±∞ or NaN
                            dst_exp = 15'h7FFF;
                            if (fp32_in[22:0] == 23'd0) begin
                                dst_mant = 64'h8000000000000000;  // ±∞
                            end else begin
                                dst_mant = {1'b1, fp32_in[22:0], 40'd0};  // NaN
                            end
                        end else begin
                            // Normalized
                            dst_exp = src_exp + 15'd16256;
                            dst_mant = {1'b1, fp32_in[22:0], 40'd0};
                        end

                        fp80_out = {dst_sign, dst_exp, dst_mant};
                        done = 1'b1;
                    end

                    //=============================================
                    // FP64 → FP80
                    //=============================================
                    MODE_FP64_TO_FP80: begin
                        // Unpack FP64
                        src_sign = fp64_in[63];
                        src_exp = {4'd0, fp64_in[62:52]};
                        src_mant = {fp64_in[51:0], 12'd0};  // Fraction only

                        dst_sign = src_sign;

                        // Handle special values
                        if (fp64_in[62:52] == 11'd0) begin
                            // Zero or denormalized
                            if (fp64_in[51:0] == 52'd0) begin
                                // ±0
                                dst_exp = 15'd0;
                                dst_mant = 64'd0;
                            end else begin
                                // Denormalized: normalize for FP80
                                shift_amount = 7'd0;
                                for (i = 51; i >= 0; i = i - 1) begin
                                    if (fp64_in[i] && shift_amount == 7'd0)
                                        shift_amount = 7'd51 - i[6:0];
                                end
                                dst_exp = 15'd16383 - 15'd1022 - {8'd0, shift_amount};
                                dst_mant = src_mant << (shift_amount + 7'd1);
                            end
                        end else if (fp64_in[62:52] == 11'd2047) begin
                            // ±∞ or NaN
                            dst_exp = 15'h7FFF;
                            if (fp64_in[51:0] == 52'd0) begin
                                dst_mant = 64'h8000000000000000;  // ±∞
                            end else begin
                                dst_mant = {1'b1, fp64_in[51:0], 11'd0};  // NaN
                            end
                        end else begin
                            // Normalized
                            dst_exp = src_exp + 15'd15360;
                            dst_mant = {1'b1, fp64_in[51:0], 11'd0};
                        end

                        fp80_out = {dst_sign, dst_exp, dst_mant};
                        done = 1'b1;
                    end

                    //=============================================
                    // FP80 → FP32
                    //=============================================
                    MODE_FP80_TO_FP32: begin
                        // Unpack FP80
                        src_sign = fp80_in[79];
                        src_exp = fp80_in[78:64];
                        src_mant = fp80_in[63:0];

                        dst_sign = src_sign;

                        // Handle special values
                        if (src_exp == 15'h7FFF) begin
                            // ±∞ or NaN
                            if (src_mant[62:0] == 63'd0 && src_mant[63] == 1'b1) begin
                                fp32_out = {dst_sign, 8'hFF, 23'd0};  // ±∞
                            end else begin
                                fp32_out = {dst_sign, 8'hFF, 1'b1, src_mant[62:41]};  // NaN
                                flag_invalid = 1'b1;
                            end
                        end else if (src_exp == 15'd0) begin
                            // ±0 or denormal
                            fp32_out = {dst_sign, 8'd0, 23'd0};
                            if (src_mant != 64'd0)
                                flag_inexact = 1'b1;
                        end else begin
                            // Normal number
                            src_exp_unbiased = {2'b00, src_exp} - 17'sd16383;

                            // Check overflow
                            if (src_exp_unbiased > 17'sd127) begin
                                fp32_out = {dst_sign, 8'hFF, 23'd0};  // ±∞
                                flag_overflow = 1'b1;
                            end else if (src_exp_unbiased < -17'sd126) begin
                                // Underflow
                                fp32_out = {dst_sign, 8'd0, 23'd0};
                                flag_underflow = 1'b1;
                                flag_inexact = 1'b1;
                            end else begin
                                // Normal range: apply rounding
                                round_up = compute_round_fp32(src_mant[39:0], rounding_mode, src_sign, src_mant[40]);

                                if (src_mant[39:0] != 40'd0)
                                    flag_inexact = 1'b1;

                                if (round_up) begin
                                    shifted_mant = {1'b1, src_mant[62:40]} + 24'd1;
                                    if (shifted_mant[24]) begin
                                        // Mantissa overflow
                                        dst_exp = (src_exp_unbiased[7:0] + 8'd127) + 8'd1;
                                        fp32_out = {dst_sign, dst_exp[7:0], shifted_mant[23:1]};
                                    end else begin
                                        dst_exp = src_exp_unbiased[7:0] + 8'd127;
                                        fp32_out = {dst_sign, dst_exp[7:0], shifted_mant[22:0]};
                                    end
                                end else begin
                                    dst_exp = src_exp_unbiased[7:0] + 8'd127;
                                    fp32_out = {dst_sign, dst_exp[7:0], src_mant[62:40]};
                                end
                            end
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // FP80 → FP64
                    //=============================================
                    MODE_FP80_TO_FP64: begin
                        // Unpack FP80
                        src_sign = fp80_in[79];
                        src_exp = fp80_in[78:64];
                        src_mant = fp80_in[63:0];

                        dst_sign = src_sign;

                        // Handle special values
                        if (src_exp == 15'h7FFF) begin
                            // ±∞ or NaN
                            if (src_mant[62:0] == 63'd0 && src_mant[63] == 1'b1) begin
                                fp64_out = {dst_sign, 11'h7FF, 52'd0};  // ±∞
                            end else begin
                                fp64_out = {dst_sign, 11'h7FF, 1'b1, src_mant[62:12]};  // NaN
                                flag_invalid = 1'b1;
                            end
                        end else if (src_exp == 15'd0) begin
                            // ±0 or denormal
                            fp64_out = {dst_sign, 11'd0, 52'd0};
                            if (src_mant != 64'd0)
                                flag_inexact = 1'b1;
                        end else begin
                            // Normal number
                            src_exp_unbiased = {2'b00, src_exp} - 17'sd16383;

                            // Check overflow
                            if (src_exp_unbiased > 17'sd1023) begin
                                fp64_out = {dst_sign, 11'h7FF, 52'd0};  // ±∞
                                flag_overflow = 1'b1;
                            end else if (src_exp_unbiased < -17'sd1022) begin
                                // Underflow
                                fp64_out = {dst_sign, 11'd0, 52'd0};
                                flag_underflow = 1'b1;
                                flag_inexact = 1'b1;
                            end else begin
                                // Normal range: apply rounding
                                round_up = compute_round_fp64(src_mant[10:0], rounding_mode, src_sign, src_mant[11]);

                                if (src_mant[10:0] != 11'd0)
                                    flag_inexact = 1'b1;

                                if (round_up) begin
                                    shifted_mant = {1'b1, src_mant[62:11]} + 53'd1;
                                    if (shifted_mant[53]) begin
                                        // Mantissa overflow
                                        dst_exp = (src_exp_unbiased[10:0] + 11'd1023) + 11'd1;
                                        fp64_out = {dst_sign, dst_exp[10:0], shifted_mant[52:1]};
                                    end else begin
                                        dst_exp = src_exp_unbiased[10:0] + 11'd1023;
                                        fp64_out = {dst_sign, dst_exp[10:0], shifted_mant[51:0]};
                                    end
                                end else begin
                                    dst_exp = src_exp_unbiased[10:0] + 11'd1023;
                                    fp64_out = {dst_sign, dst_exp[10:0], src_mant[62:11]};
                                end
                            end
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // Int16 → FP80
                    //=============================================
                    MODE_INT16_TO_FP80: begin
                        if (int16_in == 16'd0) begin
                            fp80_out = 80'd0;
                        end else begin
                            // Get sign and absolute value
                            dst_sign = int16_in[15];
                            abs_int_value = dst_sign ? (-int16_in) : int16_in;

                            // Find leading 1
                            shift_amount = 7'd0;
                            for (i = 15; i >= 0; i = i - 1) begin
                                if (abs_int_value[i] && shift_amount == 7'd0)
                                    shift_amount = 7'd15 - i[6:0];
                            end

                            // Calculate exponent
                            dst_exp = 15'd16383 + (15'd15 - {8'd0, shift_amount});

                            // Normalize mantissa
                            dst_mant = {abs_int_value[15:0], 48'd0} << shift_amount;

                            fp80_out = {dst_sign, dst_exp, dst_mant};
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // Int32 → FP80
                    //=============================================
                    MODE_INT32_TO_FP80: begin
                        if (int32_in == 32'd0) begin
                            fp80_out = 80'd0;
                        end else begin
                            // Get sign and absolute value
                            dst_sign = int32_in[31];
                            abs_int_value = dst_sign ? (-int32_in) : int32_in;

                            // Find leading 1
                            shift_amount = 7'd0;
                            for (i = 31; i >= 0; i = i - 1) begin
                                if (abs_int_value[i] && shift_amount == 7'd0)
                                    shift_amount = 7'd31 - i[6:0];
                            end

                            // Calculate exponent
                            dst_exp = 15'd16383 + (15'd31 - {8'd0, shift_amount});

                            // Normalize mantissa
                            dst_mant = {abs_int_value[31:0], 32'd0} << shift_amount;

                            fp80_out = {dst_sign, dst_exp, dst_mant};
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // FP80 → Int16
                    //=============================================
                    MODE_FP80_TO_INT16: begin
                        // Unpack FP80
                        src_sign = fp80_in[79];
                        src_exp = fp80_in[78:64];
                        src_mant = fp80_in[63:0];

                        // Handle special values
                        if (src_exp == 15'h7FFF) begin
                            // ±∞ or NaN
                            flag_invalid = 1'b1;
                            int16_out = src_sign ? 16'sh8000 : 16'sh7FFF;
                        end else if (src_exp == 15'd0) begin
                            // ±0 or denormal
                            int16_out = 16'd0;
                            if (src_mant != 64'd0)
                                flag_inexact = 1'b1;
                        end else begin
                            // Normal number
                            src_exp_unbiased = {2'b00, src_exp} - 17'sd16383;

                            if (src_exp_unbiased > 17'sd15) begin
                                // Overflow - too large for int16, set invalid (not overflow)
                                flag_invalid = 1'b1;
                                int16_out = src_sign ? 16'sh8000 : 16'sh7FFF;
                            end else if (src_exp_unbiased < -17'sd1) begin
                                // Fractional value
                                int16_out = 16'd0;
                                flag_inexact = 1'b1;
                            end else begin
                                // Convert
                                shift_amount = 7'd63 - src_exp_unbiased[6:0];
                                shifted_mant = src_mant >> shift_amount;
                                signed_int_value = shifted_mant[15:0];

                                // Check inexact
                                if (shift_amount > 7'd0 && (src_mant & ((64'd1 << shift_amount) - 64'd1)) != 64'd0) begin
                                    flag_inexact = 1'b1;
                                    round_up = compute_round_int(rounding_mode, src_sign, shift_amount > 7'd0 ? src_mant[shift_amount - 7'd1] : 1'b0);
                                    if (round_up)
                                        signed_int_value = signed_int_value + 64'd1;
                                end

                                // Apply sign
                                if (src_sign)
                                    signed_int_value = -signed_int_value;

                                // Check overflow after rounding
                                if (signed_int_value > 64'sd32767 || signed_int_value < -64'sd32768) begin
                                    flag_invalid = 1'b1;  // Set invalid for integer overflow
                                    int16_out = src_sign ? 16'sh8000 : 16'sh7FFF;
                                end else begin
                                    int16_out = signed_int_value[15:0];
                                end
                            end
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // FP80 → Int32
                    //=============================================
                    MODE_FP80_TO_INT32: begin
                        // Unpack FP80
                        src_sign = fp80_in[79];
                        src_exp = fp80_in[78:64];
                        src_mant = fp80_in[63:0];

                        // Handle special values
                        if (src_exp == 15'h7FFF) begin
                            // ±∞ or NaN
                            flag_invalid = 1'b1;
                            int32_out = src_sign ? 32'sh80000000 : 32'sh7FFFFFFF;
                        end else if (src_exp == 15'd0) begin
                            // ±0 or denormal
                            int32_out = 32'd0;
                            if (src_mant != 64'd0)
                                flag_inexact = 1'b1;
                        end else begin
                            // Normal number
                            src_exp_unbiased = {2'b00, src_exp} - 17'sd16383;

                            if (src_exp_unbiased > 17'sd31) begin
                                // Overflow - too large for int32, set invalid (not overflow)
                                flag_invalid = 1'b1;
                                int32_out = src_sign ? 32'sh80000000 : 32'sh7FFFFFFF;
                            end else if (src_exp_unbiased < -17'sd1) begin
                                // Fractional value
                                int32_out = 32'd0;
                                flag_inexact = 1'b1;
                            end else begin
                                // Convert
                                shift_amount = 7'd63 - src_exp_unbiased[6:0];
                                shifted_mant = src_mant >> shift_amount;
                                signed_int_value = shifted_mant[31:0];

                                // Check inexact
                                if (shift_amount > 7'd0 && (src_mant & ((64'd1 << shift_amount) - 64'd1)) != 64'd0) begin
                                    flag_inexact = 1'b1;
                                    round_up = compute_round_int(rounding_mode, src_sign, shift_amount > 7'd0 ? src_mant[shift_amount - 7'd1] : 1'b0);
                                    if (round_up)
                                        signed_int_value = signed_int_value + 64'd1;
                                end

                                // Apply sign
                                if (src_sign)
                                    signed_int_value = -signed_int_value;

                                // Check overflow after rounding
                                if (signed_int_value > 64'sd2147483647 || signed_int_value < -64'sd2147483648) begin
                                    flag_invalid = 1'b1;  // Set invalid for integer overflow
                                    int32_out = src_sign ? 32'sh80000000 : 32'sh7FFFFFFF;
                                end else begin
                                    int32_out = signed_int_value[31:0];
                                end
                            end
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // UInt64 → FP80
                    //=============================================
                    MODE_UINT64_TO_FP80: begin
                        if (uint64_in == 64'd0) begin
                            fp80_out = 80'd0;
                        end else begin
                            dst_sign = uint64_sign;

                            // Find leading 1
                            shift_amount = 7'd0;
                            for (i = 63; i >= 0; i = i - 1) begin
                                if (uint64_in[i] && shift_amount == 7'd0)
                                    shift_amount = 7'd63 - i[6:0];
                            end

                            // Calculate exponent
                            dst_exp = 15'd16383 + (15'd63 - {8'd0, shift_amount});

                            // Normalize mantissa
                            dst_mant = uint64_in << shift_amount;

                            fp80_out = {dst_sign, dst_exp, dst_mant};
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // FP80 → UInt64
                    //=============================================
                    MODE_FP80_TO_UINT64: begin
                        // Unpack FP80
                        src_sign = fp80_in[79];
                        src_exp = fp80_in[78:64];
                        src_mant = fp80_in[63:0];

                        uint64_sign_out = src_sign;

                        // Handle special values
                        if (src_exp == 15'h7FFF) begin
                            // ±∞ or NaN
                            flag_invalid = 1'b1;
                            uint64_out = 64'hFFFFFFFFFFFFFFFF;
                        end else if (src_exp == 15'd0) begin
                            // ±0 or denormal
                            uint64_out = 64'd0;
                            if (src_mant != 64'd0)
                                flag_inexact = 1'b1;
                        end else begin
                            // Normal number
                            src_exp_unbiased = {2'b00, src_exp} - 17'sd16383;

                            if (src_exp_unbiased > 17'sd63) begin
                                // Overflow
                                flag_overflow = 1'b1;
                                uint64_out = 64'hFFFFFFFFFFFFFFFF;
                            end else if (src_exp_unbiased < -17'sd1) begin
                                // Fractional value
                                uint64_out = 64'd0;
                                flag_inexact = 1'b1;
                            end else begin
                                // Convert
                                shift_amount = 7'd63 - src_exp_unbiased[6:0];
                                shifted_mant = src_mant >> shift_amount;
                                abs_int_value = shifted_mant;

                                // Check inexact
                                if (shift_amount > 7'd0 && (src_mant & ((64'd1 << shift_amount) - 64'd1)) != 64'd0) begin
                                    flag_inexact = 1'b1;
                                    round_up = compute_round_uint(rounding_mode, shift_amount > 7'd0 ? src_mant[shift_amount - 7'd1] : 1'b0);
                                    if (round_up) begin
                                        if (abs_int_value == 64'hFFFFFFFFFFFFFFFF)
                                            flag_overflow = 1'b1;
                                        else
                                            abs_int_value = abs_int_value + 64'd1;
                                    end
                                end

                                uint64_out = abs_int_value;
                            end
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // FP80 → Q2.62 Fixed-Point
                    //=============================================
                    MODE_FP80_TO_FIXED64: begin
                        // Unpack FP80
                        src_sign = fp80_in[79];
                        src_exp = fp80_in[78:64];
                        src_mant = fp80_in[63:0];

                        // Q2.62 format: 2 integer bits, 62 fractional bits
                        // Value = fixed_val / 2^62
                        // FP80: value = mantissa * 2^(exp - 16383 - 63)
                        // We want: fixed_val = value * 2^62
                        //        = mantissa * 2^(exp - 16383 - 63 + 62)
                        //        = mantissa * 2^(exp - 16384)

                        // Handle special values
                        if (src_exp == 15'd0) begin
                            // Zero or denormal
                            fixed64_out = 64'd0;
                        end else if (src_exp == 15'h7FFF) begin
                            // ±∞ or NaN
                            flag_invalid = 1'b1;
                            fixed64_out = 64'd0;
                        end else begin
                            // Normalized value
                            src_exp_unbiased = {2'b0, src_exp} - 17'd16384;

                            // Check for overflow (value >= 2 or <= -2)
                            if (src_exp_unbiased >= 17'sd1) begin
                                flag_overflow = 1'b1;
                                // Saturate to max/min Q2.62 value
                                if (src_sign)
                                    fixed64_out = 64'h8000000000000000;  // Most negative
                                else
                                    fixed64_out = 64'h7FFFFFFFFFFFFFFF;  // Most positive
                            end else if (src_exp_unbiased < -17'sd62) begin
                                // Underflow to zero
                                flag_underflow = 1'b1;
                                fixed64_out = 64'd0;
                            end else begin
                                // Normal conversion
                                if (src_exp_unbiased >= 0) begin
                                    // Left shift
                                    shifted_mant = src_mant << src_exp_unbiased[5:0];
                                    flag_inexact = 1'b0;
                                end else begin
                                    // Right shift
                                    shift_amount = -src_exp_unbiased[6:0];
                                    shifted_mant = src_mant >> shift_amount;
                                    // Check if bits were lost
                                    if ((src_mant & ((64'd1 << shift_amount) - 64'd1)) != 64'd0)
                                        flag_inexact = 1'b1;
                                end

                                // Check for overflow after shift (value exceeds signed 64-bit range)
                                if (!src_sign && shifted_mant >= 64'h8000000000000000) begin
                                    // Positive value >= 2.0 (MSB set means >= 2^63)
                                    flag_overflow = 1'b1;
                                    fixed64_out = 64'h7FFFFFFFFFFFFFFF;  // Saturate to max
                                end else if (src_sign && shifted_mant > 64'h8000000000000000) begin
                                    // Negative value < -2.0 (magnitude > 2^63)
                                    flag_overflow = 1'b1;
                                    fixed64_out = 64'h8000000000000000;  // Saturate to min
                                end else begin
                                    // Apply sign
                                    if (src_sign)
                                        fixed64_out = -$signed(shifted_mant);
                                    else
                                        fixed64_out = $signed(shifted_mant);
                                end
                            end
                        end
                        done = 1'b1;
                    end

                    //=============================================
                    // Q2.62 Fixed-Point → FP80
                    //=============================================
                    MODE_FIXED64_TO_FP80: begin
                        // Q2.62 format: value = fixed_val / 2^62
                        // FP80: value = mantissa * 2^(exp - 16383 - 63)

                        signed_int_value = $signed(fixed64_in);

                        if (signed_int_value == 64'sd0) begin
                            // Zero
                            fp80_out = 80'd0;
                        end else begin
                            // Extract sign
                            dst_sign = signed_int_value[63];
                            abs_int_value = dst_sign ? -signed_int_value : signed_int_value;

                            // Find leading one (normalization)
                            shift_amount = 7'd0;
                            for (i = 63; i >= 0; i = i - 1) begin
                                if (abs_int_value[i] && shift_amount == 7'd0)
                                    shift_amount = 7'd63 - i[6:0];
                            end

                            // Normalize mantissa (shift so MSB is 1)
                            dst_mant = abs_int_value << shift_amount;

                            // Compute exponent
                            // After normalization: dst_mant[63] = 1
                            // FP80 value = dst_mant * 2^(exp - 16383 - 63)
                            // We want: dst_mant * 2^(exp - 16446) = abs_int_value / 2^62
                            // => dst_mant << shift_amount = abs_int_value
                            // => (abs_int_value >> shift_amount) * 2^(exp - 16446) = abs_int_value / 2^62
                            // => 2^(exp - 16446) = 2^(-62 - shift_amount)
                            // => exp = 16384 - shift_amount
                            dst_exp = 15'd16384 - {8'd0, shift_amount};

                            fp80_out = {dst_sign, dst_exp, dst_mant};
                        end
                        done = 1'b1;
                    end

                    default: begin
                        // Invalid mode
                        done = 1'b1;
                        flag_invalid = 1'b1;
                    end
                endcase
            end else begin
                done = 1'b0;
            end
        end
    end

    //=================================================================
    // Rounding Functions
    //=================================================================

    function compute_round_fp32;
        input [39:0] discarded_bits;
        input [1:0]  rmode;
        input        sign;
        input        lsb;  // LSB of result (for round-to-even)
        begin
            compute_round_fp32 = 1'b0;
            if (discarded_bits != 40'd0) begin
                case (rmode)
                    2'b00: begin  // Round to nearest
                        if (discarded_bits[39]) begin  // Guard bit
                            if (discarded_bits[38:0] != 39'd0)
                                compute_round_fp32 = 1'b1;
                            else
                                compute_round_fp32 = lsb;  // Tie: round to even
                        end
                    end
                    2'b01: compute_round_fp32 = sign;    // Round down
                    2'b10: compute_round_fp32 = !sign;   // Round up
                    2'b11: compute_round_fp32 = 1'b0;    // Truncate
                endcase
            end
        end
    endfunction

    function compute_round_fp64;
        input [10:0] discarded_bits;
        input [1:0]  rmode;
        input        sign;
        input        lsb;
        begin
            compute_round_fp64 = 1'b0;
            if (discarded_bits != 11'd0) begin
                case (rmode)
                    2'b00: begin  // Round to nearest
                        if (discarded_bits[10]) begin  // Guard bit
                            if (discarded_bits[9:0] != 10'd0)
                                compute_round_fp64 = 1'b1;
                            else
                                compute_round_fp64 = lsb;  // Tie: round to even
                        end
                    end
                    2'b01: compute_round_fp64 = sign;
                    2'b10: compute_round_fp64 = !sign;
                    2'b11: compute_round_fp64 = 1'b0;
                endcase
            end
        end
    endfunction

    function compute_round_int;
        input [1:0]  rmode;
        input        sign;
        input        guard_bit;
        begin
            compute_round_int = 1'b0;
            case (rmode)
                2'b00: compute_round_int = guard_bit;  // Round to nearest
                2'b01: compute_round_int = sign;       // Round down
                2'b10: compute_round_int = !sign;      // Round up
                2'b11: compute_round_int = 1'b0;       // Truncate
            endcase
        end
    endfunction

    function compute_round_uint;
        input [1:0]  rmode;
        input        guard_bit;
        begin
            compute_round_uint = 1'b0;
            case (rmode)
                2'b00: compute_round_uint = guard_bit;  // Round to nearest
                2'b01: compute_round_uint = 1'b0;       // Round down
                2'b10: compute_round_uint = 1'b1;       // Round up
                2'b11: compute_round_uint = 1'b0;       // Truncate
            endcase
        end
    endfunction

endmodule
