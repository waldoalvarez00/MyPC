// Copyright 2025, Waldo Alvarez, https://pipflow.com
`timescale 1ns / 1ps

//=====================================================================
// Newton-Raphson Square Root Module (not instantiated in production build;
// SQRT is handled via microcode to save area, left as reference)
//
// Computes square root using Newton-Raphson iteration:
// x_{n+1} = 0.5 * (x_n + S/x_n)
//
// Where S is the input value and x_n converges to √S.
//
// Algorithm:
// 1. Generate initial approximation from exponent
// 2. Iterate: x_new = (x + S/x) / 2
// 3. Converge when |x_new - x| < threshold
// 4. Return result
//
// Typical convergence: 10-15 iterations for 64-bit precision
//=====================================================================

module FPU_SQRT_Newton(
    input wire clk,
    input wire reset,

    // Control
    input wire enable,

    // Input (80-bit FP)
    input wire [79:0] s_in,         // Value to take square root of

    // Output (80-bit FP)
    output reg [79:0] sqrt_out,

    output reg done,
    output reg error                // Error if s_in < 0, ±∞, or NaN
);

    //=================================================================
    // Parameters
    //=================================================================

    localparam MAX_ITERATIONS = 15;  // Maximum Newton-Raphson iterations

    //=================================================================
    // Constants
    //=================================================================

    localparam FP80_ZERO      = 80'h0000_0000000000000000;
    localparam FP80_ONE       = 80'h3FFF_8000000000000000;
    localparam FP80_HALF      = 80'h3FFE_8000000000000000;  // 0.5
    localparam FP80_TWO       = 80'h4000_8000000000000000;  // 2.0

    //=================================================================
    // State Machine
    //=================================================================

    localparam STATE_IDLE       = 4'd0;
    localparam STATE_CHECK      = 4'd1;
    localparam STATE_INIT_APPROX= 4'd2;
    localparam STATE_DIVIDE     = 4'd3;
    localparam STATE_WAIT_DIV   = 4'd4;
    localparam STATE_ADD        = 4'd5;
    localparam STATE_WAIT_ADD   = 4'd6;
    localparam STATE_MULTIPLY   = 4'd7;
    localparam STATE_WAIT_MUL   = 4'd8;
    localparam STATE_DONE       = 4'd9;

    reg [3:0] state;

    //=================================================================
    // Working Registers
    //=================================================================

    reg [79:0] s_value;         // Input value S
    reg [79:0] x_current;       // Current approximation
    reg [79:0] x_next;          // Next approximation
    reg [4:0] iteration_count;  // Iteration counter

    //=================================================================
    // Input Analysis
    //=================================================================

    wire sign_in   = s_in[79];
    wire [14:0] exp_in  = s_in[78:64];
    wire [63:0] mant_in = s_in[63:0];

    wire is_zero = (exp_in == 15'd0) && (mant_in == 64'd0);
    wire is_inf  = (exp_in == 15'h7FFF) && (mant_in[63] == 1'b1) && (mant_in[62:0] == 63'd0);
    wire is_nan  = (exp_in == 15'h7FFF) && ((mant_in[63] == 1'b0) || (mant_in[62:0] != 63'd0));
    wire is_negative = sign_in && !is_zero;

    //=================================================================
    // Arithmetic Units
    //=================================================================

    // Divide: S / x_current
    reg div_enable;
    wire [79:0] div_result;
    wire div_done;
    wire div_invalid, div_div_by_zero, div_overflow, div_underflow, div_inexact;
    reg [79:0] div_operand_a, div_operand_b;

    FPU_IEEE754_Divide div_unit (
        .clk(clk),
        .reset(reset),
        .enable(div_enable),
        .operand_a(div_operand_a),
        .operand_b(div_operand_b),
        .rounding_mode(2'b00),  // Round to nearest (default)
        .result(div_result),
        .done(div_done),
        .flag_invalid(div_invalid),
        .flag_div_by_zero(div_div_by_zero),
        .flag_overflow(div_overflow),
        .flag_underflow(div_underflow),
        .flag_inexact(div_inexact)
    );

    // Add: x_current + (S / x_current)
    reg add_enable;
    wire [79:0] add_result;
    wire add_done;
    wire add_cmp_equal, add_cmp_less, add_cmp_greater;
    wire add_invalid, add_overflow, add_underflow, add_inexact;
    reg [79:0] add_operand_a, add_operand_b;

    FPU_IEEE754_AddSub add_unit (
        .clk(clk),
        .reset(reset),
        .enable(add_enable),
        .operand_a(add_operand_a),
        .operand_b(add_operand_b),
        .subtract(1'b0),  // Addition only
        .rounding_mode(2'b00),  // Round to nearest
        .result(add_result),
        .done(add_done),
        .cmp_equal(add_cmp_equal),
        .cmp_less(add_cmp_less),
        .cmp_greater(add_cmp_greater),
        .flag_invalid(add_invalid),
        .flag_overflow(add_overflow),
        .flag_underflow(add_underflow),
        .flag_inexact(add_inexact)
    );

    // Multiply: result * 0.5
    reg mul_enable;
    wire [79:0] mul_result;
    wire mul_done;
    wire mul_invalid, mul_overflow, mul_underflow, mul_inexact;
    reg [79:0] mul_operand_a, mul_operand_b;

    FPU_IEEE754_Multiply mul_unit (
        .clk(clk),
        .reset(reset),
        .enable(mul_enable),
        .operand_a(mul_operand_a),
        .operand_b(mul_operand_b),
        .rounding_mode(2'b00),  // Round to nearest
        .result(mul_result),
        .done(mul_done),
        .flag_invalid(mul_invalid),
        .flag_overflow(mul_overflow),
        .flag_underflow(mul_underflow),
        .flag_inexact(mul_inexact)
    );

    //=================================================================
    // Initial Approximation
    //
    // Use exponent-based approximation:
    // If S = 2^E × M, then √S ≈ 2^(E/2) × √M
    // For M ∈ [1, 2), √M ∈ [1, √2), approximate as 1.0
    // So initial approximation: x₀ = 2^(E/2)
    //=================================================================

    function [79:0] initial_approximation;
        input [79:0] s;
        reg sign;
        reg [14:0] exponent;
        reg [63:0] mantissa;
        reg [14:0] sqrt_exp;
        reg [79:0] result;
        begin
            sign = s[79];
            exponent = s[78:64];
            mantissa = s[63:0];

            if (exponent == 15'd0) begin
                // Zero or denormal
                result = FP80_ZERO;
            end else begin
                // Compute √exponent
                // Subtract bias, divide by 2, add bias back
                // exp_unbiased = exponent - 16383
                // sqrt_exp = (exp_unbiased / 2) + 16383
                // = (exponent - 16383) / 2 + 16383
                // = exponent/2 + 16383/2
                // = (exponent + 16383) / 2

                sqrt_exp = (exponent + 16383) >> 1;  // Divide by 2

                // Use mantissa 1.0 (0x8000000000000000) as initial guess
                result = {1'b0, sqrt_exp, 64'h8000000000000000};
            end

            initial_approximation = result;
        end
    endfunction

    //=================================================================
    // Main State Machine
    //=================================================================

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= STATE_IDLE;
            done <= 1'b0;
            error <= 1'b0;
            sqrt_out <= FP80_ZERO;
            s_value <= FP80_ZERO;
            x_current <= FP80_ZERO;
            x_next <= FP80_ZERO;
            iteration_count <= 5'd0;
            div_enable <= 1'b0;
            add_enable <= 1'b0;
            mul_enable <= 1'b0;
        end else begin
            case (state)
                STATE_IDLE: begin
                    done <= 1'b0;
                    error <= 1'b0;
                    div_enable <= 1'b0;
                    add_enable <= 1'b0;
                    mul_enable <= 1'b0;

                    if (enable) begin
                        s_value <= s_in;
                        state <= STATE_CHECK;
                    end
                end

                STATE_CHECK: begin
                    // Check for special cases
                    if (is_negative) begin
                        // Error: square root of negative number
                        error <= 1'b1;
                        state <= STATE_DONE;
                    end else if (is_zero) begin
                        // √0 = 0
                        sqrt_out <= FP80_ZERO;
                        state <= STATE_DONE;
                    end else if (is_inf) begin
                        // √∞ = ∞
                        sqrt_out <= s_value;
                        state <= STATE_DONE;
                    end else if (is_nan) begin
                        // √NaN = NaN
                        sqrt_out <= s_value;
                        state <= STATE_DONE;
                    end else begin
                        // Normal case: proceed with Newton-Raphson
                        state <= STATE_INIT_APPROX;
                    end
                end

                STATE_INIT_APPROX: begin
                    // Generate initial approximation
                    x_current <= initial_approximation(s_value);
                    iteration_count <= 5'd0;
                    state <= STATE_DIVIDE;
                end

                STATE_DIVIDE: begin
                    // Compute S / x_current
                    div_operand_a <= s_value;
                    div_operand_b <= x_current;
                    div_enable <= 1'b1;
                    state <= STATE_WAIT_DIV;
                end

                STATE_WAIT_DIV: begin
                    div_enable <= 1'b0;
                    if (div_done) begin
                        // Store S/x for next step
                        state <= STATE_ADD;
                    end
                end

                STATE_ADD: begin
                    // Compute x_current + (S / x_current)
                    add_operand_a <= x_current;
                    add_operand_b <= div_result;
                    add_enable <= 1'b1;
                    state <= STATE_WAIT_ADD;
                end

                STATE_WAIT_ADD: begin
                    add_enable <= 1'b0;
                    if (add_done) begin
                        // Store sum for next step
                        state <= STATE_MULTIPLY;
                    end
                end

                STATE_MULTIPLY: begin
                    // Compute 0.5 * (x_current + S/x_current)
                    mul_operand_a <= add_result;
                    mul_operand_b <= FP80_HALF;
                    mul_enable <= 1'b1;
                    state <= STATE_WAIT_MUL;
                end

                STATE_WAIT_MUL: begin
                    mul_enable <= 1'b0;
                    if (mul_done) begin
                        x_next <= mul_result;

                        // Check iteration count
                        iteration_count <= iteration_count + 1;
                        if (iteration_count >= MAX_ITERATIONS - 1) begin
                            // Max iterations reached, return result
                            sqrt_out <= mul_result;
                            state <= STATE_DONE;
                        end else begin
                            // Continue iterating
                            x_current <= mul_result;
                            state <= STATE_DIVIDE;
                        end
                    end
                end

                STATE_DONE: begin
                    done <= 1'b1;
                    if (~enable) begin
                        state <= STATE_IDLE;
                    end
                end

                default: state <= STATE_IDLE;
            endcase
        end
    end

endmodule


//=====================================================================
// IMPLEMENTATION NOTES
//=====================================================================
//
// This is a FUNCTIONAL Newton-Raphson square root with placeholder arithmetic.
//
// TO COMPLETE INTEGRATION:
//
// 1. Connect Real Divide Unit:
//    FPU_IEEE754_Divide div_unit (
//        .clk(clk),
//        .reset(reset),
//        .enable(div_enable),
//        .operand_a(div_operand_a),
//        .operand_b(div_operand_b),
//        .result(div_result),
//        .done(div_done),
//        ...
//    );
//
// 2. Connect Real Add Unit:
//    FPU_IEEE754_AddSub add_unit (
//        .clk(clk),
//        .reset(reset),
//        .enable(add_enable),
//        .operand_a(add_operand_a),
//        .operand_b(add_operand_b),
//        .subtract(1'b0),
//        .result(add_result),
//        .done(add_done),
//        ...
//    );
//
// 3. Connect Real Multiply Unit:
//    FPU_IEEE754_Multiply mul_unit (
//        .clk(clk),
//        .reset(reset),
//        .enable(mul_enable),
//        .operand_a(mul_operand_a),
//        .operand_b(mul_operand_b),
//        .result(mul_result),
//        .done(mul_done),
//        ...
//    );
//
// 4. Add Convergence Check:
//    Current version uses fixed iteration count (15 iterations).
//    Enhancement: Check if |x_next - x_current| < threshold
//    to terminate early when converged.
//
// 5. Optimize Initial Approximation:
//    Current: Uses exponent-based approximation
//    Enhancement: Use lookup table for better initial guess
//    to reduce iteration count.
//
// PERFORMANCE:
// - Typical: 10-12 iterations for convergence
// - Each iteration: 1 divide (~60 cycles) + 1 add (~10 cycles) + 1 multiply (~25 cycles)
//   ≈ 95 cycles per iteration
// - Total: ~950-1140 cycles (comparable to real 8087 FSQRT at ~180-200 cycles)
// - Can be optimized with better initial approximation
//
// TESTING STRATEGY:
// 1. Test perfect squares: √4 = 2, √9 = 3, √16 = 4
// 2. Test powers of 2: √2, √8, √32
// 3. Test small values: √0.25 = 0.5, √0.0625 = 0.25
// 4. Compare against Python math.sqrt()
// 5. Verify error cases: √(-1) should set error flag
//=====================================================================


//=====================================================================
// NEWTON-RAPHSON CONVERGENCE ANALYSIS
//=====================================================================
//
// Newton-Raphson for √S:
//   f(x) = x² - S
//   f'(x) = 2x
//   x_{n+1} = x_n - f(x_n)/f'(x_n)
//          = x_n - (x_n² - S)/(2x_n)
//          = (2x_n² - x_n² + S)/(2x_n)
//          = (x_n² + S)/(2x_n)
//          = (x_n + S/x_n)/2
//
// Convergence rate: Quadratic (doubles precision each iteration)
//
// Error analysis:
//   e_n = x_n - √S (error at iteration n)
//   e_{n+1} ≈ e_n²/(2√S)
//
// Starting with 8-bit accuracy (from exponent approximation):
//   Iteration 1: 16-bit accuracy
//   Iteration 2: 32-bit accuracy
//   Iteration 3: 64-bit accuracy (sufficient for FP80 mantissa)
//   Iterations 4-5: Refinement to eliminate rounding errors
//
// Therefore, 10-15 iterations provides more than sufficient precision
// for 80-bit extended precision floating point.
//=====================================================================
