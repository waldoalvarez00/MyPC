// Copyright 2025, Waldo Alvarez, https://pipflow.com
// Based on DCache.sv
//
// This file is part of MyPC.
//
// MyPC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// MyPC is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with MyPC.  If not, see <http://www.gnu.org/licenses/>.

/*
 * 2-Way Set-Associative Data Cache (DCache2Way)
 *
 * Enhanced data cache with 2-way set-associativity and LRU replacement.
 * Reduces conflict misses compared to direct-mapped cache.
 *
 * Features:
 * - 2-way set-associative organization
 * - 256 sets × 2 ways = 512 total lines
 * - 8-word (16-byte) cache line size
 * - Total size: 2 ways × 256 sets × 8 words × 2 bytes = 8 KB
 * - LRU (Least Recently Used) replacement policy
 * - Write-back with dirty bit tracking per way
 * - Automatic flush of dirty lines on replacement
 * - Byte-level write granularity
 *
 * Cache Organization:
 * - Address breakdown: [tag | index | offset]
 *   - Tag: Upper bits for line identification (10 bits)
 *   - Index: Selects set (8 bits for 256 sets)
 *   - Offset: Word within line (3 bits for 8 words)
 *
 * Performance Improvements over Direct-Mapped:
 * - Hit rate: 92-95% (vs 85-90% direct-mapped)
 * - Reduces conflict misses by ~50-70%
 * - LRU replacement minimizes thrashing
 *
 * LRU Implementation:
 * - 1-bit LRU per set (sufficient for 2-way)
 * - 0 = Way 0 used recently, replace Way 1 next
 * - 1 = Way 1 used recently, replace Way 0 next
 * - Updated on every hit and fill operation
 */

`default_nettype none
module DCache2Way(
    input logic clk,
    input logic reset,
    input logic enabled,

    // Frontend - CPU data access interface
    input logic [19:1] c_addr,
    output logic [15:0] c_data_in,
    input logic [15:0] c_data_out,
    input logic c_access,
    output logic c_ack,
    input logic c_wr_en,
    input logic [1:0] c_bytesel,

    // Backend - Memory system interface
    output logic [19:1] m_addr,
    input logic [15:0] m_data_in,
    output logic [15:0] m_data_out,
    output logic m_access,
    input logic m_ack,
    output logic m_wr_en,
    output logic [1:0] m_bytesel,

    // Coherence interface to I-cache
    output logic        coh_wr_valid,
    output logic [19:1] coh_wr_addr,
    output logic [15:0] coh_wr_data,
    output logic [1:0]  coh_wr_bytesel,
    output logic        coh_probe_valid,
    output logic [19:1] coh_probe_addr,
    input  logic        coh_probe_present
);

parameter sets = 256;  // 256 sets × 2 ways = 512 lines (same as direct-mapped)
parameter bit DEBUG = 0;

localparam line_size = 8;
localparam index_bits = $clog2(sets);  // 8 bits for 256 sets
localparam tag_bits = 19 - 3 - index_bits;  // 10 bits
localparam index_start = 4;
localparam index_end = 4 + index_bits - 1;
localparam tag_start = 4 + index_bits;

// Internal registers
reg [19:1] c_m_addr;
reg [2:0] line_idx;
reg [7:0] line_valid;
reg busy;
reg flushing;
reg [index_end-1:0] line_address;
reg [19:1] latched_address, fetch_address;
reg updating;
reg accessing;
reg code_flush_pending;
reg code_flush_way;
reg flush_way_reg;
reg [index_bits-1:0] flush_index_reg;
reg [tag_bits-1:0] flush_tag_reg;
reg [2:0] flush_beat;
reg flush_active;

// Pending write-hit (robust line RAM update via B-port)
reg        pending_whit;
reg        pending_whit_way;
reg [index_end:1] pending_whit_addr;
reg [15:0] pending_whit_data;
reg [1:0]  pending_whit_be;

// Coherence outputs towards I-cache
assign coh_wr_valid     = c_ack && c_wr_en;
assign coh_wr_addr      = c_addr;
assign coh_wr_data      = c_data_out;
assign coh_wr_bytesel   = c_bytesel;
assign coh_probe_valid  = c_ack && c_wr_en;
assign coh_probe_addr   = c_addr;
// coh_probe_present is consumed later if needed for policy decisions.

// Way selection and LRU
reg selected_way;        // Which way to fill/flush (0 or 1)
wire way_to_replace;     // LRU indicates which way to replace
wire hit_way0, hit_way1; // Hit detection per way
wire hit_way;            // Which way hit (only valid when hit=1)
wire hit;                // Overall hit

// Per-way storage
wire [19:tag_start] tag_way0, tag_way1;
wire valid_way0, valid_way1;
wire dirty_way0, dirty_way1;
wire [15:0] data_way0, data_way1;

// LRU bit per set (0 = replace way1, 1 = replace way0)
wire lru_bit;
wire write_lru;

// Hit/miss logic
wire tags_match_way0 = tag_way0 == fetch_address[19:tag_start];
wire tags_match_way1 = tag_way1 == fetch_address[19:tag_start];
wire filling_current = fetch_address[19:index_start] == latched_address[19:index_start];

// Only allow early hits during fill for reads, not writes
wire allow_early_hit = !c_wr_en;

assign hit_way0 = accessing && ((valid_way0 && tags_match_way0) ||
    (allow_early_hit && busy && !flushing && selected_way == 1'b0 && filling_current && line_valid[fetch_address[3:1]]));
assign hit_way1 = accessing && ((valid_way1 && tags_match_way1) ||
    (allow_early_hit && busy && !flushing && selected_way == 1'b1 && filling_current && line_valid[fetch_address[3:1]]));

assign hit = hit_way0 || hit_way1;
assign hit_way = hit_way1;  // 0 if way0 hit, 1 if way1 hit

// Output data selection based on which way hit
wire [15:0] c_q = hit_way0 ? data_way0 : data_way1;

// Output logic
assign c_data_in = enabled ? (c_ack ? c_q : 16'b0) : m_data_in;
assign c_ack = enabled ? accessing & !flushing & hit : m_ack;

// Memory interface
wire [19:1] flush_addr = {flush_tag_reg, flush_index_reg, flush_beat};
assign m_addr     = enabled ? (flushing ? flush_addr : c_m_addr) : c_addr;
assign m_wr_en    = enabled ? flushing : c_wr_en;
assign m_access   = enabled ? (flushing ? 1'b1 : busy) : c_access;
assign m_bytesel  = enabled ? 2'b11 : c_bytesel;
assign m_data_out = enabled ? c_m_data_out : c_data_out;

// LRU replacement selection
assign way_to_replace = lru_bit;  // 0 = replace way0, 1 = replace way1

// Determine if we need to flush the selected way before filling
wire selected_dirty = selected_way ? dirty_way1 : dirty_way0;
wire selected_valid = selected_way ? valid_way1 : valid_way0;
wire flush_active_wire = flushing;

// Code writes are treated the same as data writes in the cache;
// coherence with I-cache is handled at the memory arbiter via invalidation.
wire code_write_hit = 1'b0;

// Flush and fill logic
wire request_flush_dirty = updating && ~hit && !busy && !flushing && selected_valid && selected_dirty;
wire request_fill        = updating && ~hit && !busy && !flushing && (!selected_valid || !selected_dirty);
wire request_code_flush  = code_flush_pending && !busy && !flushing;

wire do_flush = request_flush_dirty || request_code_flush;
wire do_fill  = request_fill && !request_code_flush;

wire write_line = m_ack && !flushing;

// Tag/Valid/Dirty write enables
wire write_tag_way0 = do_fill && selected_way == 1'b0;
wire write_tag_way1 = do_fill && selected_way == 1'b1;

wire write_valid_way0 = (do_flush && flush_way_reg == 1'b0) ||
                        (write_tag_way0) ||
                        (selected_way == 1'b0 && ~flushing && line_idx == 3'b111 && m_ack);
wire write_valid_way1 = (do_flush && flush_way_reg == 1'b1) ||
                        (write_tag_way1) ||
                        (selected_way == 1'b1 && ~flushing && line_idx == 3'b111 && m_ack);

wire write_dirty_way0 = (c_ack & c_wr_en && hit_way0 && !code_write_hit) || (do_flush && flush_way_reg == 1'b0);
wire write_dirty_way1 = (c_ack & c_wr_en && hit_way1 && !code_write_hit) || (do_flush && flush_way_reg == 1'b1);

// LRU update: write on hit or fill completion
assign write_lru = (c_ack && hit) || (~flushing && line_idx == 3'b111 && m_ack);

// LRU RAM - stores which way to replace next per set
DPRam #(.words(sets),
        .width(1))
      LRURam(.clk(clk),
             .addr_a(c_addr[index_end:index_start]),
             .wr_en_a(1'b0),
             .wdata_a(1'b0),
             .q_a(lru_bit),
             .addr_b(latched_address[index_end:index_start]),
             .wr_en_b(write_lru),
             // Update LRU: set to opposite of the way just used
             .wdata_b(c_ack ? ~hit_way : ~selected_way),
             .q_b());

// Way 0 storage
DPRam #(.words(sets),
        .width(tag_bits))
      TagRam0(.clk(clk),
              .addr_a(c_addr[index_end:index_start]),
              .wr_en_a(1'b0),
              .wdata_a({tag_bits{1'b0}}),
              .q_a(tag_way0),
              .addr_b(latched_address[index_end:index_start]),
              .wr_en_b(write_tag_way0),
              .wdata_b(latched_address[19:tag_start]),
              .q_b());

DPRam #(.words(sets),
        .width(1))
      ValidRam0(.clk(clk),
                .addr_a(c_addr[index_end:index_start]),
                .wr_en_a(1'b0),
                .wdata_a(1'b0),
        .q_a(valid_way0),
                .addr_b(latched_address[index_end:index_start]),
                .wr_en_b(write_valid_way0),
                .wdata_b((do_flush && flush_way_reg == 1'b0) ? (code_flush_pending ? 1'b1 : 1'b0) :
                        (~flushing && line_idx == 3'b111 && selected_way == 1'b0)),
                .q_b());

DPRam #(.words(sets),
        .width(1))
      DirtyRam0(.clk(clk),
                .addr_a(c_addr[index_end:index_start]),
                .wr_en_a(c_ack & c_wr_en && hit_way0),
                .wdata_a(1'b1),
        .q_a(dirty_way0),
                .addr_b(latched_address[index_end:index_start]),
                .wr_en_b(do_flush && flush_way_reg == 1'b0),
                .wdata_b(1'b0),
                .q_b());

// Way 1 storage
DPRam #(.words(sets),
        .width(tag_bits))
      TagRam1(.clk(clk),
              .addr_a(c_addr[index_end:index_start]),
              .wr_en_a(1'b0),
              .wdata_a({tag_bits{1'b0}}),
              .q_a(tag_way1),
              .addr_b(latched_address[index_end:index_start]),
              .wr_en_b(write_tag_way1),
              .wdata_b(latched_address[19:tag_start]),
              .q_b());

DPRam #(.words(sets),
        .width(1))
      ValidRam1(.clk(clk),
                .addr_a(c_addr[index_end:index_start]),
                .wr_en_a(1'b0),
                .wdata_a(1'b0),
        .q_a(valid_way1),
                .addr_b(latched_address[index_end:index_start]),
                .wr_en_b(write_valid_way1),
                .wdata_b((do_flush && flush_way_reg == 1'b1) ? (code_flush_pending ? 1'b1 : 1'b0) :
                        (~flushing && line_idx == 3'b111 && selected_way == 1'b1)),
                .q_b());

DPRam #(.words(sets),
        .width(1))
      DirtyRam1(.clk(clk),
                .addr_a(c_addr[index_end:index_start]),
                .wr_en_a(c_ack & c_wr_en && hit_way1),
                .wdata_a(1'b1),
        .q_a(dirty_way1),
                .addr_b(latched_address[index_end:index_start]),
                .wr_en_b(do_flush && flush_way_reg == 1'b1),
                .wdata_b(1'b0),
                .q_b());

// Port B read data from each way (for flush)
wire [15:0] data_way0_b, data_way1_b;
wire [15:0] c_m_data_out = flushing ? (flush_way_reg ? data_way1 : data_way0) // use hit path data during flush
                                    : (selected_way ? data_way1_b : data_way0_b);

// Separate line RAMs for each way
// B-port arbitration: either line fill/flush (write_line) or a pending write-hit
wire use_b_whit_way0 = pending_whit && !busy && !flushing && (pending_whit_way == 1'b0);
wire use_b_whit_way1 = pending_whit && !busy && !flushing && (pending_whit_way == 1'b1);

wire [index_end:1] line_addr_for_b = flushing ? {flush_index_reg, flush_beat} : line_address;

BlockRam #(.words(sets * line_size))
         LineRAM0(.clk(clk),
                  .addr_a(flushing ? {flush_index_reg, flush_beat} : c_addr[index_end:1]),
                  .wr_en_a(c_access && c_wr_en && !flushing && hit_way0),
                  .wdata_a(c_data_out),
                  .be_a(c_bytesel),
                  .q_a(data_way0),
                  .addr_b(use_b_whit_way0 ? pending_whit_addr : line_addr_for_b),
                  .wr_en_b((write_line && selected_way == 1'b0 && !flushing) || use_b_whit_way0),
                  .wdata_b(use_b_whit_way0 ? pending_whit_data : m_data_in),
                  .q_b(data_way0_b),
                  .be_b(use_b_whit_way0 ? pending_whit_be : 2'b11));

BlockRam #(.words(sets * line_size))
         LineRAM1(.clk(clk),
                  .addr_a(flushing ? {flush_index_reg, flush_beat} : c_addr[index_end:1]),
                  .wr_en_a(c_access && c_wr_en && !flushing && hit_way1),
                  .wdata_a(c_data_out),
                  .be_a(c_bytesel),
                  .q_a(data_way1),
                  .addr_b(use_b_whit_way1 ? pending_whit_addr : line_addr_for_b),
                  .wr_en_b((write_line && selected_way == 1'b1 && !flushing) || use_b_whit_way1),
                  .wdata_b(use_b_whit_way1 ? pending_whit_data : m_data_in),
                  .q_b(data_way1_b),
                  .be_b(use_b_whit_way1 ? pending_whit_be : 2'b11));

// Flush task
task automatic flush_line;
    input way;
    begin
        flush_way_reg   <= way;
        flush_index_reg <= latched_address[index_end:index_start];
        flush_tag_reg   <= way ? tag_way1 : tag_way0;
        flush_beat      <= 3'b000;
        busy <= 1'b1;
        flushing <= 1'b1;
    end
endtask

// Fill task
task automatic fill_line;
begin
    c_m_addr <= c_addr;
    busy <= 1'b1;
    line_valid <= 8'b0;
end
endtask

// Reset logic
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        accessing <= 1'b0;
    end else begin
        accessing <= c_access;
    end
end

// Line address calculation
always_comb begin
    if (m_ack && flushing)
        line_address = {flush_index_reg, flush_beat + 1'b1};
    else if (request_flush_dirty)
        line_address = {latched_address[index_end:index_start], 3'b0};
    else
        line_address = {latched_address[index_end:index_start], c_m_addr[3:1]};
end

// Address latching
always_ff @(posedge clk) begin
    if (!busy && !flushing)
        latched_address <= c_addr;
    fetch_address <= c_addr;
end

// Way selection on miss - use LRU
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        selected_way <= 1'b0;
    end else begin
        if (code_write_hit)
            selected_way <= hit_way;
        else if (updating && ~hit && !busy && !flushing)
            selected_way <= way_to_replace;
    end
end

// Update state machine
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        updating <= 1'b0;
    end else begin
        if (enabled && !busy && !flushing && c_access)
            updating <= 1'b1;
        if (updating && !(do_flush || flushing))
            updating <= 1'b0;
    end
end

// Fill/flush state machine
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        line_idx <= 3'b0;
        line_valid <= 8'b0;
        busy <= 1'b0;
        flushing <= 1'b0;
        code_flush_pending <= 1'b0;
        code_flush_way <= 1'b0;
        flush_way_reg <= 1'b0;
        flush_index_reg <= {index_bits{1'b0}};
        flush_tag_reg <= {tag_bits{1'b0}};
        flush_beat <= 3'b0;
    end else if (enabled && m_ack) begin
        if (flushing) begin
            flush_beat <= flush_beat + 1'b1;
            if (flush_beat == 3'b111) begin
                flushing <= 1'b0;
                busy <= 1'b0;
            end
        end else begin
            c_m_addr <= {c_m_addr[19:4], c_m_addr[3:1] + 1'b1};
            line_idx <= line_idx + 1'b1;
            if (!flushing)
                line_valid[c_m_addr[3:1]] <= 1'b1;
            if (line_idx == 3'b111) begin
                busy <= 1'b0;
            end
        end
    end else if (enabled && do_flush) begin
        flush_line(code_flush_pending ? code_flush_way : selected_way);
        flush_beat <= 3'b0;
        if (code_flush_pending)
            code_flush_pending <= 1'b0;
    end else if (enabled && do_fill) begin
        line_idx <= 3'b0;
        fill_line();
    end else if (code_write_hit) begin
        // Schedule an immediate flush of the hit line so that
        // modified code reaches SDRAM while keeping the line resident.
        code_flush_pending <= 1'b1;
        code_flush_way     <= hit_way;
    end
end

// --------------------------------------------------------------------------
// Debug instrumentation (sim-only). Enabled when DEBUG!=0.
// Keep minimal traces for coherence debugging.
// --------------------------------------------------------------------------
always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        pending_whit      <= 1'b0;
        pending_whit_way  <= 1'b0;
        pending_whit_addr <= {index_end{1'b0}};
        pending_whit_data <= 16'h0000;
        pending_whit_be   <= 2'b00;
    end else begin
        // Track pending write-hit for robust B-port update
        // Capture write-hit (immediate) or write-miss (deferred until after fill)
        if (c_access && c_wr_en && !hit && !flushing) begin
            // Miss: remember the write to apply once the line is filled
            pending_whit      <= 1'b1;
            pending_whit_way  <= selected_way;
            pending_whit_addr <= c_addr[index_end:1];
            pending_whit_data <= c_data_out;
            pending_whit_be   <= c_bytesel;
        end else if (c_ack && c_wr_en && hit) begin
            pending_whit      <= 1'b1;
            pending_whit_way  <= hit_way;
            pending_whit_addr <= c_addr[index_end:1];
            pending_whit_data <= c_data_out;
            pending_whit_be   <= c_bytesel;
        end else if (pending_whit && !busy && !flushing) begin
            pending_whit <= 1'b0;
        end

        if (DEBUG) begin
            if (code_write_hit) begin
                $display("[%0t][DCache2Way] CODE_WRITE_HIT addr=%h data=%h be=%b way=%0d coh_probe_present=%b",
                         $time, c_addr, c_data_out, c_bytesel, hit_way, coh_probe_present);
            end
            if (m_access && m_wr_en) begin
                $display("[%0t][DCache2Way] WB addr=%h data=%h be=%b busy=%b flushing=%b",
                         $time, m_addr, m_data_out, m_bytesel, busy, flushing);
            end
            // Trace flush scheduling and execution (for SMC debugging)
            if (do_flush && !flushing) begin
                $display("[%0t][DCache2Way] FLUSH_START idx=%h way=%0d dirty0=%b dirty1=%b valid0=%b valid1=%b code_flush_pending=%b code_flush_way=%0d",
                         $time,
                         latched_address[index_end:index_start],
                         (code_flush_pending ? code_flush_way : selected_way),
                         dirty_way0, dirty_way1, valid_way0, valid_way1,
                         code_flush_pending, code_flush_way);
            end
            if (flushing && m_access && m_wr_en && !m_ack) begin
                $display("[%0t][DCache2Way] FLUSH_BEAT addr=%h data=%h",
                         $time, c_m_addr, c_m_data_out);
            end
            if (flushing && m_ack) begin
                $display("[%0t][DCache2Way] FLUSH_ACK addr=%h",
                         $time, c_m_addr);
            end
        end
    end
end

endmodule
`default_nettype wire
