`timescale 1ns / 1ps

//=====================================================================
// Test for Control Instructions: FINIT, FLDCW, FSTCW, FSTSW
//
// Tests:
// - FINIT: Initialize FPU (reset stack, control word, status word)
// - FLDCW: Load control word from memory
// - FSTCW: Store control word to memory
// - FSTSW: Store status word to memory
//=====================================================================

module tb_control_instructions;

    // Clock and reset
    reg clk;
    reg reset;

    // FPU Core signals
    reg [7:0]   instruction;
    reg [2:0]   stack_index;
    reg         execute;
    wire        ready;
    wire        error;
    reg [79:0]  data_in;
    wire [79:0] data_out;
    reg [31:0]  int_data_in;
    wire [31:0] int_data_out;

    // Memory operand format
    reg         has_memory_op;
    reg [1:0]   operand_size;
    reg         is_integer;
    reg         is_bcd;

    // Control/Status interface
    reg [15:0]  control_in;
    reg         control_write;
    wire [15:0] status_out;
    wire [15:0] control_out;
    wire [15:0] tag_word_out;

    // Test tracking
    integer test_count, pass_count, fail_count;

    //=================================================================
    // FPU Core Instantiation
    //=================================================================

    FPU_Core fpu (
        .clk(clk),
        .reset(reset),
        .instruction(instruction),
        .stack_index(stack_index),
        .execute(execute),
        .ready(ready),
        .error(error),
        .data_in(data_in),
        .data_out(data_out),
        .int_data_in(int_data_in),
        .int_data_out(int_data_out),
        .has_memory_op(has_memory_op),
        .operand_size(operand_size),
        .is_integer(is_integer),
        .is_bcd(is_bcd),
        .control_in(control_in),
        .control_write(control_write),
        .status_out(status_out),
        .control_out(control_out),
        .tag_word_out(tag_word_out)
    );

    //=================================================================
    // Clock Generation
    //=================================================================

    always begin
        #5 clk = ~clk;
    end

    //=================================================================
    // Test Tasks
    //=================================================================

    // Execute FPU instruction
    task execute_instruction;
        input [7:0] op;
        input [79:0] data;
        begin
            @(posedge clk);
            instruction <= op;
            stack_index <= 3'd0;
            data_in <= data;
            int_data_in <= 32'd0;
            has_memory_op <= 1'b0;
            operand_size <= 2'd0;
            is_integer <= 1'b0;
            is_bcd <= 1'b0;
            control_in <= 16'd0;
            control_write <= 1'b0;
            execute <= 1'b1;
            @(posedge clk);
            execute <= 1'b0;

            // Wait for ready
            wait(ready);
            @(posedge clk);
            // Extra cycles to allow register outputs to settle
            @(posedge clk);
            @(posedge clk);
        end
    endtask

    // Test FINIT instruction
    task test_finit;
        input [255:0] test_name;
        begin
            test_count = test_count + 1;
            $display("[Test %0d] %s", test_count, test_name);

            // Execute FINIT
            execute_instruction(8'hF0, 80'd0);

            // Check results
            if (tag_word_out == 16'hFFFF &&  // All tags empty (0b11 per register)
                control_out == 16'h037F &&  // Default control word
                status_out[5:0] == 6'd0) begin  // Exception flags cleared
                $display("  PASS: tag_word=0x%h, control_word=0x%h, status=0x%h",
                         tag_word_out, control_out, status_out);
                pass_count = pass_count + 1;
            end else begin
                $display("  FAIL: tag_word=0x%h (expected 0xFFFF)",
                         tag_word_out);
                $display("        control_word=0x%h (expected 0x037F), status_word=0x%h",
                         control_out, status_out);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Test FLDCW instruction
    task test_fldcw;
        input [255:0] test_name;
        input [15:0] control_value;
        begin
            test_count = test_count + 1;
            $display("[Test %0d] %s", test_count, test_name);

            // Execute FLDCW with control word in data_in[15:0]
            execute_instruction(8'hF1, {64'd0, control_value});

            // Wait one more cycle for control_out to update
            @(posedge clk);

            // Check that control word was loaded
            if (control_out == control_value) begin
                $display("  PASS: control_word=0x%h", control_out);
                pass_count = pass_count + 1;
            end else begin
                $display("  FAIL: control_word=0x%h (expected 0x%h)",
                         control_out, control_value);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Test FSTCW instruction
    task test_fstcw;
        input [255:0] test_name;
        input [15:0] expected_control;
        begin
            test_count = test_count + 1;
            $display("[Test %0d] %s", test_count, test_name);

            // Execute FSTCW
            execute_instruction(8'hF2, 80'd0);

            // Check that control word was stored to outputs
            if (int_data_out[15:0] == expected_control &&
                data_out[15:0] == expected_control) begin
                $display("  PASS: int_data_out=0x%h, data_out[15:0]=0x%h",
                         int_data_out[15:0], data_out[15:0]);
                pass_count = pass_count + 1;
            end else begin
                $display("  FAIL: int_data_out=0x%h, data_out[15:0]=0x%h (expected 0x%h)",
                         int_data_out[15:0], data_out[15:0], expected_control);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Test FSTSW instruction
    task test_fstsw;
        input [255:0] test_name;
        begin
            test_count = test_count + 1;
            $display("[Test %0d] %s", test_count, test_name);

            // Execute FSTSW
            execute_instruction(8'hF3, 80'd0);

            // Check that status word was stored to outputs
            if (int_data_out[15:0] == status_out &&
                data_out[15:0] == status_out) begin
                $display("  PASS: int_data_out=0x%h, data_out[15:0]=0x%h, status=0x%h",
                         int_data_out[15:0], data_out[15:0], status_out);
                pass_count = pass_count + 1;
            end else begin
                $display("  FAIL: int_data_out=0x%h, data_out[15:0]=0x%h, status=0x%h",
                         int_data_out[15:0], data_out[15:0], status_out);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Test FNINIT instruction (no-wait version)
    task test_finit_nowait;
        input [255:0] test_name;
        begin
            test_count = test_count + 1;
            $display("[Test %0d] %s", test_count, test_name);

            // Execute FNINIT (opcode 0xF6)
            execute_instruction(8'hF6, 80'd0);

            // Check results (same as FINIT)
            if (tag_word_out == 16'hFFFF &&  // All tags empty (0b11 per register)
                control_out == 16'h037F &&  // Default control word
                status_out[5:0] == 6'd0) begin  // Exception flags cleared
                $display("  PASS: tag_word=0x%h, control_word=0x%h, status=0x%h",
                         tag_word_out, control_out, status_out);
                pass_count = pass_count + 1;
            end else begin
                $display("  FAIL: tag_word=0x%h (expected 0xFFFF)",
                         tag_word_out);
                $display("        control_word=0x%h (expected 0x037F), status_word=0x%h",
                         control_out, status_out);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Test FNSTCW instruction (no-wait version)
    task test_fstcw_nowait;
        input [255:0] test_name;
        input [15:0] expected_control;
        begin
            test_count = test_count + 1;
            $display("[Test %0d] %s", test_count, test_name);

            // Execute FNSTCW (opcode 0xF7)
            execute_instruction(8'hF7, 80'd0);

            // Check that control word was stored to outputs
            if (int_data_out[15:0] == expected_control &&
                data_out[15:0] == expected_control) begin
                $display("  PASS: int_data_out=0x%h, data_out[15:0]=0x%h",
                         int_data_out[15:0], data_out[15:0]);
                pass_count = pass_count + 1;
            end else begin
                $display("  FAIL: int_data_out=0x%h, data_out[15:0]=0x%h (expected 0x%h)",
                         int_data_out[15:0], data_out[15:0], expected_control);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Test FNSTSW instruction (no-wait version)
    task test_fstsw_nowait;
        input [255:0] test_name;
        begin
            test_count = test_count + 1;
            $display("[Test %0d] %s", test_count, test_name);

            // Execute FNSTSW (opcode 0xF8)
            execute_instruction(8'hF8, 80'd0);

            // Check that status word was stored to outputs
            if (int_data_out[15:0] == status_out &&
                data_out[15:0] == status_out) begin
                $display("  PASS: int_data_out=0x%h, data_out[15:0]=0x%h, status=0x%h",
                         int_data_out[15:0], data_out[15:0], status_out);
                pass_count = pass_count + 1;
            end else begin
                $display("  FAIL: int_data_out=0x%h, data_out[15:0]=0x%h, status=0x%h",
                         int_data_out[15:0], data_out[15:0], status_out);
                fail_count = fail_count + 1;
            end
        end
    endtask

    //=================================================================
    // Main Test Sequence
    //=================================================================

    initial begin
        // Initialize
        clk = 0;
        reset = 1;
        instruction = 8'd0;
        stack_index = 3'd0;
        execute = 0;
        data_in = 80'd0;
        int_data_in = 32'd0;
        has_memory_op = 1'b0;
        operand_size = 2'd0;
        is_integer = 1'b0;
        is_bcd = 1'b0;
        control_in = 16'd0;
        control_write = 1'b0;

        test_count = 0;
        pass_count = 0;
        fail_count = 0;

        // Reset
        #20;
        reset = 0;
        #20;

        $display("\nControl Instructions Test Suite");
        $display("==================================================\n");

        // ===========================
        // FINIT Tests
        // ===========================
        $display("Testing FINIT (Initialize FPU)");
        $display("--------------------------------------------------");

        // Test 1: FINIT should reset everything
        test_finit("FINIT - Initialize FPU");

        $display("");

        // ===========================
        // FLDCW Tests
        // ===========================
        $display("Testing FLDCW (Load Control Word)");
        $display("--------------------------------------------------");

        // Test 2: Load default control word
        test_fldcw("FLDCW - Load default (0x037F)", 16'h037F);

        // Test 3: Load control word with different rounding mode
        test_fldcw("FLDCW - Round down (0x077F)", 16'h077F);

        // Test 4: Load control word with different precision
        test_fldcw("FLDCW - Single precision (0x007F)", 16'h007F);

        // Test 5: Load control word with exceptions unmasked
        test_fldcw("FLDCW - Unmask all exceptions (0x0300)", 16'h0300);

        $display("");

        // ===========================
        // FSTCW Tests
        // ===========================
        $display("Testing FSTCW (Store Control Word)");
        $display("--------------------------------------------------");

        // Test 6: Store current control word (should be 0x0300 from test 5)
        test_fstcw("FSTCW - Store control word", 16'h0300);

        // Test 7: Load new value and store it
        test_fldcw("FLDCW - Load 0x0FFF", 16'h0FFF);
        test_fstcw("FSTCW - Store 0x0FFF", 16'h0FFF);

        $display("");

        // ===========================
        // FSTSW Tests
        // ===========================
        $display("Testing FSTSW (Store Status Word)");
        $display("--------------------------------------------------");

        // Test 8: Store status word
        test_fstsw("FSTSW - Store status word");

        // Test 9: Store status word after FINIT
        execute_instruction(8'hF0, 80'd0);  // FINIT
        test_fstsw("FSTSW - Store after FINIT");

        $display("");

        // ===========================
        // No-Wait Instruction Tests
        // ===========================
        $display("Testing No-Wait Versions (FNINIT, FNSTCW, FNSTSW)");
        $display("--------------------------------------------------");

        // Test 11: FNINIT (no-wait version of FINIT)
        test_finit_nowait("FNINIT - Initialize FPU (no-wait)");

        // Test 12: FNSTCW (no-wait version of FSTCW)
        execute_instruction(8'hF1, {64'd0, 16'h0BCD});  // FLDCW first
        @(posedge clk);
        test_fstcw_nowait("FNSTCW - Store control word (no-wait)", 16'h0BCD);

        // Test 13: FNSTSW (no-wait version of FSTSW)
        test_fstsw_nowait("FNSTSW - Store status word (no-wait)");

        $display("");

        // ===========================
        // Integration Tests
        // ===========================
        $display("Testing Integration Scenarios");
        $display("--------------------------------------------------");

        // Test 14: FINIT + FLDCW + FSTCW sequence
        test_count = test_count + 1;
        $display("[Test %0d] FINIT + FLDCW + FSTCW sequence", test_count);

        execute_instruction(8'hF0, 80'd0);  // FINIT
        execute_instruction(8'hF1, {64'd0, 16'h0A5A});  // FLDCW
        execute_instruction(8'hF2, 80'd0);  // FSTCW

        if (control_out == 16'h0A5A && int_data_out[15:0] == 16'h0A5A) begin
            $display("  PASS: Control word sequence works correctly");
            pass_count = pass_count + 1;
        end else begin
            $display("  FAIL: control_word=0x%h, stored=0x%h (expected 0x0A5A)",
                     control_out, int_data_out[15:0]);
            fail_count = fail_count + 1;
        end

        // Test 15: Verify FINIT resets control word
        test_count = test_count + 1;
        $display("[Test %0d] FINIT resets control word to 0x037F", test_count);

        execute_instruction(8'hF1, {64'd0, 16'hFFFF});  // FLDCW with all bits set
        execute_instruction(8'hF0, 80'd0);  // FINIT

        // Wait for control word to update
        @(posedge clk);

        if (control_out == 16'h037F) begin
            $display("  PASS: FINIT correctly resets control word");
            pass_count = pass_count + 1;
        end else begin
            $display("  FAIL: control_word=0x%h (expected 0x037F)", control_out);
            fail_count = fail_count + 1;
        end

        $display("");

        // ===========================
        // Summary
        // ===========================
        $display("==================================================");
        $display("Test Summary");
        $display("==================================================");
        $display("Total tests:  %0d", test_count);
        $display("Passed:       %0d", pass_count);
        $display("Failed:       %0d", fail_count);
        $display("");

        if (fail_count == 0) begin
            $display("*** ALL TESTS PASSED ***");
        end else begin
            $display("*** %0d TEST(S) FAILED ***", fail_count);
        end
        $display("");

        $finish;
    end

endmodule
