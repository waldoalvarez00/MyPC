`timescale 1ns/1ps

module floppy_tb;

    // Clock and reset
    logic clk;
    logic reset;

    // DMA interface
    logic dma_req;
    logic dma_ack;
    logic dma_tc;
    logic [7:0] dma_readdata;
    logic [7:0] dma_writedata;

    // IRQ
    logic irq;

    // I/O interface
    logic [2:0] io_address;
    logic io_read;
    logic [7:0] io_readdata;
    logic io_write;
    logic [7:0] io_writedata;
    logic bus_ack;

    // Media management (stubbed)
    logic [3:0] mgmt_address;
    logic mgmt_fddn;
    logic mgmt_write;
    logic [15:0] mgmt_writedata;
    logic mgmt_read;
    logic [15:0] mgmt_readdata;
    logic fdd0_inserted;

    // Other
    logic [1:0] wp;
    logic [27:0] clock_rate;
    logic [1:0] request;

    // Test tracking
    integer test_count = 0;
    integer pass_count = 0;
    integer fail_count = 0;

    // Test variables (Icarus-compatible - declared at module level)
    logic [7:0] dor_val;
    logic [7:0] msr_val;
    logic [7:0] dir_val;

    // Clock generation: 50 MHz (20ns period)
    parameter CLK_PERIOD = 20;
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end

    // DUT instantiation
    floppy dut (
        .clk(clk),
        .reset(reset),
        .dma_req(dma_req),
        .dma_ack(dma_ack),
        .dma_tc(dma_tc),
        .dma_readdata(dma_readdata),
        .dma_writedata(dma_writedata),
        .irq(irq),
        .io_address(io_address),
        .io_read(io_read),
        .io_readdata(io_readdata),
        .io_write(io_write),
        .io_writedata(io_writedata),
        .bus_ack(bus_ack),
        .fdd0_inserted(fdd0_inserted),
        .mgmt_address(mgmt_address),
        .mgmt_fddn(mgmt_fddn),
        .mgmt_write(mgmt_write),
        .mgmt_writedata(mgmt_writedata),
        .mgmt_read(mgmt_read),
        .mgmt_readdata(mgmt_readdata),
        .wp(wp),
        .clock_rate(clock_rate),
        .request(request)
    );

    // Test result checking task
    task automatic check_result(
        input string test_name,
        input logic [7:0] expected,
        input logic [7:0] actual
    );
        test_count++;
        if (expected === actual) begin
            $display("[PASS] %s: Expected 0x%02h, Got 0x%02h", test_name, expected, actual);
            pass_count++;
        end else begin
            $display("[FAIL] %s: Expected 0x%02h, Got 0x%02h", test_name, expected, actual);
            fail_count++;
        end
    endtask

    // I/O write task
    task automatic io_write_reg(
        input logic [2:0] addr,
        input logic [7:0] data
    );
        io_address = addr;
        io_writedata = data;
        io_write = 1'b1;
        io_read = 1'b0;
        @(posedge clk);
        wait (bus_ack);
        @(posedge clk);
        io_write = 1'b0;
        @(posedge clk);
    endtask

    // I/O read task
    task automatic io_read_reg(
        input logic [2:0] addr,
        output logic [7:0] data
    );
        io_address = addr;
        io_write = 1'b0;
        io_read = 1'b1;
        @(posedge clk);
        wait (bus_ack);
        @(posedge clk);
        data = io_readdata;
        io_read = 1'b0;
        @(posedge clk);
    endtask

    // Main test sequence
    initial begin
        // Initialize
        $display("================================================");
        $display("Floppy Disk Controller Testbench");
        $display("================================================\n");

        reset = 1;
        dma_ack = 0;
        dma_tc = 0;
        dma_readdata = 8'h00;
        io_address = 3'h0;
        io_read = 0;
        io_write = 0;
        io_writedata = 8'h00;
        mgmt_address = 4'h0;
        mgmt_fddn = 0;
        mgmt_write = 0;
        mgmt_writedata = 16'h0000;
        mgmt_read = 0;
        wp = 2'b00;
        clock_rate = 28'd50_000_000;

        // Wait for reset
        repeat (10) @(posedge clk);
        reset = 0;
        repeat (5) @(posedge clk);

        $display("Test 1: Digital Output Register (DOR) - Port 0x3F2");
        $display("---------------------------------------------------");

        // Test 1a: Write DOR - Enable controller, select drive 0, motors off
        io_write_reg(3'h2, 8'b0000_0100);  // DMA=0, RESET=1, DRV_SEL=0, MOTA=0, MOTB=0
        #(CLK_PERIOD * 5);

        // Test 1b: Read DOR back
        io_read_reg(3'h2, dor_val);
        check_result("DOR Write/Read", 8'b0000_0100, dor_val);

        $display("\nTest 2: Main Status Register (MSR) - Port 0x3F4");
        $display("---------------------------------------------------");

        // Test 2a: Read MSR - should show RQM=1 (ready for command)
        io_read_reg(3'h4, msr_val);
        $display("MSR Initial State: 0x%02h (RQM=%b, DIO=%b, BUSY=%b)",
                 msr_val, msr_val[7], msr_val[6], msr_val[4]);

        if (msr_val[7] == 1'b1) begin
            $display("[PASS] MSR shows ready for command (RQM=1)");
            pass_count++;
        end else begin
            $display("[FAIL] MSR should show ready (RQM=1), got RQM=%b", msr_val[7]);
            fail_count++;
        end
        test_count++;

        $display("\nTest 3: SPECIFY Command (0x03)");
        $display("---------------------------------------------------");

        // Test 3a: Send SPECIFY command (set step rate, head load/unload times)
        // Command format: 03h, [SRT:HUT], [HLT:ND]
        // SRT=4ms, HUT=8ms, HLT=16ms, ND=0 (DMA mode)
        io_write_reg(3'h5, 8'h03);        // SPECIFY command
        #(CLK_PERIOD * 5);
        io_write_reg(3'h5, 8'h48);        // SRT=4, HUT=8
        #(CLK_PERIOD * 5);
        io_write_reg(3'h5, 8'h20);        // HLT=16ms, ND=0 (DMA mode)
        #(CLK_PERIOD * 10);

        // Test 3b: Verify command completed (RQM should be 1, BUSY should be 0)
        io_read_reg(3'h4, msr_val);
        if (msr_val[7] == 1'b1 && msr_val[4] == 1'b0) begin
            $display("[PASS] SPECIFY command completed successfully");
            pass_count++;
        end else begin
            $display("[FAIL] SPECIFY command did not complete properly");
            fail_count++;
        end
        test_count++;

        $display("\nTest 4: VERSION Command (0x10)");
        $display("---------------------------------------------------");

        // Test 4a: Send VERSION command
        io_write_reg(3'h5, 8'h10);        // VERSION command
        #(CLK_PERIOD * 10);

        // Test 4b: Read version from FIFO (should return 0x90 for enhanced controller)
        io_read_reg(3'h4, msr_val);
        $display("MSR after VERSION: 0x%02h (RQM=%b, DIO=%b, BUSY=%b)",
                 msr_val, msr_val[7], msr_val[6], msr_val[4]);

        if (msr_val[6] == 1'b1) begin  // DIO=1 means result ready
            logic [7:0] version;
            io_read_reg(3'h5, version);
            check_result("VERSION", 8'h90, version);
        end else begin
            $display("[FAIL] No result available after VERSION command");
            fail_count++;
            test_count++;
        end

        $display("\nTest 5: Digital Input Register (DIR) - Port 0x3F7");
        $display("---------------------------------------------------");

        // Test 5a: Read DIR - bit 7 is disk change signal
        io_read_reg(3'h7, dir_val);
        $display("DIR Value: 0x%02h (DSKCHG=%b)", dir_val, dir_val[7]);

        // Disk change should be set (no media inserted)
        if (dir_val[7] == 1'b1) begin
            $display("[PASS] DIR shows disk change (no media)");
            pass_count++;
        end else begin
            $display("[FAIL] DIR should show disk change");
            fail_count++;
        end
        test_count++;

        $display("\nTest 6: SENSE INTERRUPT STATUS Command (0x08)");
        $display("---------------------------------------------------");

        // Test 6a: Send SENSE INTERRUPT STATUS
        io_write_reg(3'h5, 8'h08);
        #(CLK_PERIOD * 10);

        // Test 6b: Read result bytes
        io_read_reg(3'h4, msr_val);
        if (msr_val[6] == 1'b1) begin  // DIO=1
            logic [7:0] st0, pcn;
            io_read_reg(3'h5, st0);
            #(CLK_PERIOD * 5);
            io_read_reg(3'h5, pcn);
            $display("SENSE INT result: ST0=0x%02h, PCN=0x%02h", st0, pcn);
            $display("[PASS] SENSE INTERRUPT STATUS executed");
            pass_count++;
        end else begin
            $display("[FAIL] No result from SENSE INTERRUPT STATUS");
            fail_count++;
        end
        test_count++;

        $display("\nTest 7: Motor Control via DOR");
        $display("---------------------------------------------------");

        // Test 7a: Enable motor for drive 0
        io_write_reg(3'h2, 8'b0001_0100);  // DMA=0, RESET=1, DRV_SEL=0, MOTA=1
        #(CLK_PERIOD * 5);

        // Test 7b: Read back DOR
        io_read_reg(3'h2, dor_val);
        check_result("Motor Enable", 8'b0001_0100, dor_val);

        // Test 7c: Disable motor
        io_write_reg(3'h2, 8'b0000_0100);  // Motors off
        #(CLK_PERIOD * 5);

        $display("\nTest 8: Invalid Command Test");
        $display("---------------------------------------------------");

        // Test 8a: Send invalid command (should return 0x80 in result)
        io_write_reg(3'h5, 8'hFF);  // Invalid command
        #(CLK_PERIOD * 10);

        // Test 8b: Check for invalid command response
        io_read_reg(3'h4, msr_val);
        if (msr_val[6] == 1'b1) begin
            logic [7:0] result;
            io_read_reg(3'h5, result);
            check_result("Invalid Command Response", 8'h80, result);
        end

        // Test Summary
        $display("\n================================================");
        $display("Test Summary");
        $display("================================================");
        $display("Total Tests: %0d", test_count);
        $display("Passed:      %0d", pass_count);
        $display("Failed:      %0d", fail_count);
        $display("Success Rate: %0d%%", (pass_count * 100) / test_count);
        $display("================================================\n");

        if (fail_count == 0)
            $display("ALL TESTS PASSED!");
        else
            $display("SOME TESTS FAILED!");

        $finish;
    end

    // Timeout watchdog
    initial begin
        #100000;  // 100 microseconds
        $display("\n[ERROR] Test timeout!");
        $display("Test may be stuck. Aborting...\n");
        $finish;
    end

    // Waveform dump
    initial begin
        $dumpfile("floppy_tb.vcd");
        $dumpvars(0, floppy_tb);
    end

endmodule
