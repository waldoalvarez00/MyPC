//
// Dual-Port RAM Module (Verilog replacement for dpram.vhd)
//
// True dual-port RAM with independent or shared clocks
//
// Copyright (c) 2024 - MIT License
//

module dpram #(
    parameter addr_width = 8,
    parameter data_width = 8
) (
    // Single clock (always use this for simulation - dual clocks not supported)
    input                       clock,
    // Dual clocks (unused in this simulation stub - clock is always used)
    input                       clock_a,
    input                       clock_b,

    // Port A
    input  [addr_width-1:0]     address_a,
    input  [data_width-1:0]     data_a,
    input                       wren_a,
    output reg [data_width-1:0] q_a,

    // Port B
    input  [addr_width-1:0]     address_b,
    input  [data_width-1:0]     data_b,
    input                       wren_b,
    output reg [data_width-1:0] q_b
);

    // For simulation, always use the single 'clock' input
    // The clock_a/clock_b inputs are ignored (they're just compatibility ports)
    wire clka = clock;
    wire clkb = clock;

    // Memory array - initialize to zeros (not random X values)
    // verilator lint_off UNUSEDSIGNAL
    (* ram_init_file = "UNUSED" *)  // Prevent Verilator from randomizing
    reg [data_width-1:0] mem [0:(2**addr_width)-1] /* verilator public */;
    // verilator lint_on UNUSEDSIGNAL

    // Initialize memory to zeros for simulation
    // verilator lint_off BLKSEQ
    integer i;
    initial begin
        for (i = 0; i < (2**addr_width); i = i + 1) begin
            mem[i] = {data_width{1'b0}};
        end
    end
    // verilator lint_on BLKSEQ

    // Port A
    always @(posedge clka) begin
        if (wren_a) begin
            mem[address_a] <= data_a;
        end
        q_a <= mem[address_a];
    end

    // Port B
    always @(posedge clkb) begin
        if (wren_b) begin
            mem[address_b] <= data_b;
        end
        q_b <= mem[address_b];
    end

endmodule

//
// Dual-Port RAM with different widths (dpram_dif)
// Supports both single-clock and dual-clock interfaces
//
module dpram_dif #(
    parameter addr_width_a = 12,
    parameter data_width_a = 8,
    parameter addr_width_b = 11,
    parameter data_width_b = 16,
    parameter init_file = ""
) (
    // Single clock (always use this for simulation - dual clocks not supported)
    input                         clock,
    // Dual clocks (unused in this simulation stub - clock is always used)
    input                         clock_a,
    input                         clock_b,

    // Port A
    input  [addr_width_a-1:0]     address_a,
    input  [data_width_a-1:0]     data_a,
    input                         wren_a,
    output reg [data_width_a-1:0] q_a,

    // Port B
    input  [addr_width_b-1:0]     address_b,
    input  [data_width_b-1:0]     data_b,
    input                         wren_b,
    output reg [data_width_b-1:0] q_b
);

    // For simulation, always use the single 'clock' input
    // The clock_a/clock_b inputs are ignored (they're just compatibility ports)
    wire clka = clock;
    wire clkb = clock;

    // Use the larger address width for memory
    localparam mem_size = (2**addr_width_a > 2**addr_width_b) ? 2**addr_width_a : 2**addr_width_b;

    // Memory array (using 8-bit granularity)
    reg [7:0] mem [0:mem_size-1];

    // Initialize memory from file if specified
    initial begin
        if (init_file != "") begin
            $readmemh(init_file, mem);
        end
    end

    // Port A (8-bit access)
    always @(posedge clka) begin
        if (wren_a) begin
            mem[address_a] <= data_a;
        end
        q_a <= mem[address_a];
    end

    // Port B (16-bit access, assumes little-endian)
    always @(posedge clkb) begin
        if (wren_b) begin
            mem[{address_b, 1'b0}]     <= data_b[7:0];
            mem[{address_b, 1'b1}]     <= data_b[15:8];
        end
        q_b <= {mem[{address_b, 1'b1}], mem[{address_b, 1'b0}]};
    end

endmodule
