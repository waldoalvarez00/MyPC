// ================================================================
// Harvard Arbiter Timing Debug Test
// Verifies ACK timing with detailed cycle-by-cycle output
// ================================================================

`timescale 1ns/1ps

module arbiter_timing_debug;

    logic clk, reset;
    logic [19:1] icache_m_addr, dcache_m_addr;
    logic [15:0] icache_m_data_in, dcache_m_data_in;
    logic [15:0] dcache_m_data_out;
    logic icache_m_access, dcache_m_access;
    logic icache_m_ack, dcache_m_ack;
    logic dcache_m_wr_en;
    logic [1:0] dcache_m_bytesel;

    logic [19:1] mem_m_addr;
    logic [15:0] mem_m_data_in, mem_m_data_out;
    logic mem_m_access, mem_m_ack, mem_m_wr_en;
    logic [1:0] mem_m_bytesel;

    // DUT
    HarvardArbiter dut (.*);

    // Clock: 50 MHz
    initial begin
        clk = 0;
        forever #10 clk = ~clk;
    end

    // Memory model - 1 cycle latency
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            mem_m_ack <= 1'b0;
            mem_m_data_in <= 16'b0;
        end else begin
            mem_m_ack <= mem_m_access;
            if (mem_m_access && !mem_m_wr_en)
                mem_m_data_in <= {8'hAA, mem_m_addr[15:8]};
        end
    end

    // Cycle counter
    int cycle;
    always_ff @(posedge clk or posedge reset)
        if (reset) cycle <= 0;
        else cycle <= cycle + 1;

    // Test
    initial begin
        $display("================================================================");
        $display("Harvard Arbiter Timing Debug");
        $display("================================================================\n");

        // Initialize
        reset = 1;
        icache_m_addr = 0;
        icache_m_access = 0;
        dcache_m_addr = 0;
        dcache_m_access = 0;
        dcache_m_wr_en = 0;
        dcache_m_data_out = 0;
        dcache_m_bytesel = 2'b11;

        repeat(3) @(posedge clk);
        reset = 0;
        repeat(2) @(posedge clk);

        $display("--- Test: Single I-cache Request Timing ---\n");
        $display("Cycle | icache | state        | grant_i | mem     | mem   | icache");
        $display("      | access |              |         | access  | ack   | ack");
        $display("------|--------|--------------|---------|---------|-------|-------");

        // Start request
        icache_m_addr = 19'h12345;
        icache_m_access = 1;

        // Monitor for 10 cycles
        repeat(10) begin
            @(posedge clk);
            #1;  // Let signals settle
            $display(" %2d   |   %b    | %12s |    %b    |    %b    |   %b   |   %b",
                cycle,
                icache_m_access,
                dut.state.name(),
                dut.grant_icache,
                mem_m_access,
                mem_m_ack,
                icache_m_ack);
        end

        $display("\nAnalysis:");
        $display("- Request starts at cycle 0");
        $display("- State transitions to SERVING_ICACHE at cycle 1");
        $display("- mem_m_access goes high at cycle 1");
        $display("- mem_m_ack goes high at cycle 2 (1 cycle memory latency)");
        $display("- icache_m_ack goes high at cycle 3 (1 cycle arbiter ACK register)");
        $display("\nConclusion: Total latency = 3 cycles from request to ACK");

        $finish;
    end

endmodule
