/**
 * tb_cpu_fpu_integrated.v
 *
 * Comprehensive Testbench for CPU+FPU Integrated System
 *
 * Tests complete system integration:
 * - CPU executing ESC instructions
 * - Memory-mapped FPU communication
 * - FPU instruction processing
 * - BUSY signal synchronization
 * - End-to-end instruction execution
 *
 * Date: 2025-11-10
 */

`timescale 1ns / 1ps

module tb_cpu_fpu_integrated;

    //=================================================================
    // Test Infrastructure
    //=================================================================

    reg clk;
    reg reset;

    // CPU Instruction Input
    reg [7:0] cpu_instruction_opcode;
    reg [7:0] cpu_instruction_modrm;
    reg cpu_instruction_valid;
    wire cpu_instruction_ack;

    // System Memory Interface
    wire [19:0] sys_mem_addr;
    reg [15:0] sys_mem_data_in;
    wire [15:0] sys_mem_data_out;
    wire sys_mem_access;
    reg sys_mem_ack;
    wire sys_mem_wr_en;
    wire [1:0] sys_mem_bytesel;

    // System Status
    wire system_busy;
    wire fpu_interrupt;
    wire [2:0] cpu_state;
    wire [15:0] fpu_status_out;

    // Test control
    integer test_num;
    integer pass_count;
    integer fail_count;
    reg [255:0] test_name;

    //=================================================================
    // Simulated Memory
    //=================================================================

    reg [15:0] memory [0:65535];
    integer i;

    // Memory simulation with realistic timing
    reg [19:0] last_mem_addr;
    reg mem_was_accessed;

    always @(posedge clk) begin
        if (reset) begin
            sys_mem_ack <= 1'b0;
            mem_was_accessed <= 1'b0;
            last_mem_addr <= 20'h00000;
        end else begin
            if (sys_mem_access) begin
                // New address or first access
                if (sys_mem_addr != last_mem_addr || !mem_was_accessed) begin
                    sys_mem_ack <= 1'b1;
                    last_mem_addr <= sys_mem_addr;
                    mem_was_accessed <= 1'b1;

                    if (!sys_mem_wr_en) begin
                        // Read from memory
                        sys_mem_data_in <= memory[sys_mem_addr[15:1]];
                    end else begin
                        // Write to memory
                        memory[sys_mem_addr[15:1]] <= sys_mem_data_out;
                    end
                end else begin
                    sys_mem_ack <= 1'b0;
                end
            end else begin
                sys_mem_ack <= 1'b0;
                mem_was_accessed <= 1'b0;
            end
        end
    end

    //=================================================================
    // DUT Instantiation
    //=================================================================

    CPU_FPU_Integrated_System dut (
        .clk(clk),
        .reset(reset),
        .cpu_instruction_opcode(cpu_instruction_opcode),
        .cpu_instruction_modrm(cpu_instruction_modrm),
        .cpu_instruction_valid(cpu_instruction_valid),
        .cpu_instruction_ack(cpu_instruction_ack),
        .sys_mem_addr(sys_mem_addr),
        .sys_mem_data_in(sys_mem_data_in),
        .sys_mem_data_out(sys_mem_data_out),
        .sys_mem_access(sys_mem_access),
        .sys_mem_ack(sys_mem_ack),
        .sys_mem_wr_en(sys_mem_wr_en),
        .sys_mem_bytesel(sys_mem_bytesel),
        .system_busy(system_busy),
        .fpu_interrupt(fpu_interrupt),
        .cpu_state(cpu_state),
        .fpu_status_out(fpu_status_out)
    );

    //=================================================================
    // Clock Generation
    //=================================================================

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    //=================================================================
    // Test Helper Tasks
    //=================================================================

    task start_test;
        input [255:0] name;
        begin
            test_num = test_num + 1;
            test_name = name;
            $display("\n========================================");
            $display("Test %0d: %0s", test_num, name);
            $display("========================================");
        end
    endtask

    task end_test;
        input pass;
        begin
            if (pass) begin
                $display("[PASS] Test %0d: %0s", test_num, test_name);
                pass_count = pass_count + 1;
            end else begin
                $display("[FAIL] Test %0d: %0s", test_num, test_name);
                fail_count = fail_count + 1;
            end
        end
    endtask

    task reset_system;
        begin
            reset = 1;
            cpu_instruction_opcode = 8'h00;
            cpu_instruction_modrm = 8'h00;
            cpu_instruction_valid = 0;

            @(posedge clk);
            @(posedge clk);
            reset = 0;
            @(posedge clk);
        end
    endtask

    task send_instruction;
        input [7:0] opcode;
        input [7:0] modrm;
        begin
            cpu_instruction_opcode = opcode;
            cpu_instruction_modrm = modrm;
            cpu_instruction_valid = 1;
            @(posedge clk);
            #1;
            cpu_instruction_valid = 0;
        end
    endtask

    task wait_instruction_complete;
        integer timeout;
        reg completed;
        begin
            completed = 0;
            timeout = 0;
            while (!completed && timeout < 200) begin
                @(posedge clk);
                if (cpu_instruction_ack) begin
                    completed = 1;
                end
                timeout = timeout + 1;
            end

            if (timeout >= 200) begin
                $display("ERROR: Instruction timeout");
            end
        end
    endtask

    task load_memory_dword;
        input [19:0] addr;
        input [31:0] data;
        begin
            memory[addr[15:1]]     = data[15:0];
            memory[addr[15:1] + 1] = data[31:16];
        end
    endtask

    //=================================================================
    // Test Execution
    //=================================================================

    initial begin
        $display("\n");
        $display("==================================================");
        $display("CPU+FPU Integrated System Test Suite");
        $display("==================================================");

        test_num = 0;
        pass_count = 0;
        fail_count = 0;

        // Initialize memory
        for (i = 0; i < 65536; i = i + 1) begin
            memory[i] = 16'h0000;
        end

        //-------------------------------------------------------------
        // Test Category 1: Basic ESC Instruction Recognition
        //-------------------------------------------------------------

        start_test("ESC D8 instruction recognition");
        reset_system();
        send_instruction(8'hD8, 8'hC1);  // FADD ST, ST(1)
        wait_instruction_complete();
        end_test(1'b1);  // If we got here, instruction completed

        start_test("ESC D9 instruction recognition");
        reset_system();
        send_instruction(8'hD9, 8'hC0);  // FLD ST(0)
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("ESC DA instruction recognition");
        reset_system();
        send_instruction(8'hDA, 8'hC2);  // FCMOVB ST, ST(2)
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("ESC DB instruction recognition");
        reset_system();
        send_instruction(8'hDB, 8'hE3);  // FINIT
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("ESC DC instruction recognition");
        reset_system();
        send_instruction(8'hDC, 8'hC8);  // FMUL ST, ST(0)
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("ESC DD instruction recognition");
        reset_system();
        send_instruction(8'hDD, 8'hD0);  // FST ST(0)
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("ESC DE instruction recognition");
        reset_system();
        send_instruction(8'hDE, 8'hD9);  // FCOMPP
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("ESC DF instruction recognition");
        reset_system();
        send_instruction(8'hDF, 8'hE0);  // FSTSW AX
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        //-------------------------------------------------------------
        // Test Category 2: Non-ESC Instructions
        //-------------------------------------------------------------

        start_test("Non-ESC instruction (MOV)");
        reset_system();
        send_instruction(8'h89, 8'hC0);  // MOV AX, AX
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("Non-ESC instruction (ADD)");
        reset_system();
        send_instruction(8'h01, 8'hC0);  // ADD AX, AX
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        //-------------------------------------------------------------
        // Test Category 3: ESC with Memory Operands
        //-------------------------------------------------------------

        start_test("FLD dword from memory");
        reset_system();
        load_memory_dword(20'h01000, 32'h12345678);
        send_instruction(8'hD9, 8'h06);  // FLD dword ptr [mem]
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("FADD dword from memory");
        reset_system();
        load_memory_dword(20'h01000, 32'hABCDEF01);
        send_instruction(8'hD8, 8'h06);  // FADD dword ptr [mem]
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("FST dword to memory");
        reset_system();
        send_instruction(8'hD9, 8'h16);  // FST dword ptr [mem]
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        //-------------------------------------------------------------
        // Test Category 4: Back-to-Back ESC Instructions
        //-------------------------------------------------------------

        start_test("Back-to-back ESC instructions");
        reset_system();
        send_instruction(8'hD8, 8'hC1);  // FADD
        wait_instruction_complete();
        @(posedge clk);
        send_instruction(8'hD8, 8'hCA);  // FMUL
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("Three consecutive ESC instructions");
        reset_system();
        send_instruction(8'hD9, 8'hC0);  // FLD
        wait_instruction_complete();
        @(posedge clk);
        send_instruction(8'hD8, 8'hC1);  // FADD
        wait_instruction_complete();
        @(posedge clk);
        send_instruction(8'hDD, 8'hD8);  // FSTP
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        //-------------------------------------------------------------
        // Test Category 5: System State Verification
        //-------------------------------------------------------------

        start_test("System returns to idle after instruction");
        reset_system();
        send_instruction(8'hD8, 8'hC1);
        wait_instruction_complete();
        @(posedge clk);
        @(posedge clk);
        end_test(cpu_state === 3'd0);  // CPU_STATE_IDLE

        start_test("System busy during instruction processing");
        reset_system();
        send_instruction(8'hD8, 8'hC1);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        end_test(system_busy === 1'b1 || cpu_instruction_ack === 1'b1);

        //-------------------------------------------------------------
        // Test Category 6: Mixed ESC and Non-ESC Instructions
        //-------------------------------------------------------------

        start_test("ESC followed by non-ESC");
        reset_system();
        send_instruction(8'hD8, 8'hC1);  // FADD (ESC)
        wait_instruction_complete();
        @(posedge clk);
        send_instruction(8'h90, 8'h00);  // NOP (non-ESC)
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        start_test("Non-ESC followed by ESC");
        reset_system();
        send_instruction(8'h90, 8'h00);  // NOP (non-ESC)
        wait_instruction_complete();
        @(posedge clk);
        send_instruction(8'hD8, 8'hC1);  // FADD (ESC)
        wait_instruction_complete();
        @(posedge clk);
        end_test(1'b1);  // Instruction completed

        //-------------------------------------------------------------
        // Test Category 7: All ESC Opcodes Coverage
        //-------------------------------------------------------------

        start_test("ESC coverage - D8");
        reset_system();
        send_instruction(8'hD8, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        start_test("ESC coverage - D9");
        reset_system();
        send_instruction(8'hD9, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        start_test("ESC coverage - DA");
        reset_system();
        send_instruction(8'hDA, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        start_test("ESC coverage - DB");
        reset_system();
        send_instruction(8'hDB, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        start_test("ESC coverage - DC");
        reset_system();
        send_instruction(8'hDC, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        start_test("ESC coverage - DD");
        reset_system();
        send_instruction(8'hDD, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        start_test("ESC coverage - DE");
        reset_system();
        send_instruction(8'hDE, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        start_test("ESC coverage - DF");
        reset_system();
        send_instruction(8'hDF, 8'hC0);
        wait_instruction_complete();
        end_test(1'b1);  // Instruction completed

        //-------------------------------------------------------------
        // Test Results Summary
        //-------------------------------------------------------------

        $display("\n");
        $display("==================================================");
        $display("Test Suite Complete");
        $display("==================================================");
        $display("Total Tests:  %0d", test_num);
        $display("Passed:       %0d", pass_count);
        $display("Failed:       %0d", fail_count);
        $display("Pass Rate:    %0d%%", (pass_count * 100) / test_num);
        $display("==================================================");

        if (fail_count == 0) begin
            $display("\n*** ALL TESTS PASSED ***\n");
        end else begin
            $display("\n*** SOME TESTS FAILED ***\n");
        end

        $finish;
    end

    //=================================================================
    // Timeout Watchdog
    //=================================================================

    initial begin
        #2000000;  // 2ms timeout
        $display("\n*** ERROR: Test timeout ***\n");
        $finish;
    end

    //=================================================================
    // Waveform Dump
    //=================================================================

    initial begin
        $dumpfile("tb_cpu_fpu_integrated.vcd");
        $dumpvars(0, tb_cpu_fpu_integrated);
    end

endmodule
