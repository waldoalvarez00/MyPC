// Copyright 2025, Waldo Alvarez, https://pipflow.com
`timescale 1ns / 1ps

//=====================================================================
// Arctangent Lookup Table for CORDIC
//
// This ROM contains 64 entries of atan(2^-i) values in 80-bit
// IEEE 754 extended precision format.
//
// Used by CORDIC algorithms for computing trigonometric functions:
// - sin/cos (rotation mode)
// - atan (vectoring mode)
// - tan (rotation mode + division)
//
// Format: atan(2^-index) where index ∈ [0, 63]
//
// Auto-generated by generate_atan_table.py
//=====================================================================

module FPU_Atan_Table(
    input wire [5:0] index,        // Index (0-63)
    output reg [79:0] atan_value   // atan(2^-index) in FP80 format
);

    // Arctangent lookup table
    always @(*) begin
        case (index)
            6'd 0: atan_value = 80'h3FFE_C90FDAA22168C000; // atan(2^- 0) = 0.78539816339744827900 rad (45.00000°)
            6'd 1: atan_value = 80'h3FFD_ED63382B0DDA7800; // atan(2^- 1) = 0.46364760900080609352 rad (26.56505°)
            6'd 2: atan_value = 80'h3FFC_FADBAFC96406E800; // atan(2^- 2) = 0.24497866312686414347 rad (14.03624°)
            6'd 3: atan_value = 80'h3FFB_FEADD4D5617B7000; // atan(2^- 3) = 0.12435499454676143816 rad ( 7.12502°)
            6'd 4: atan_value = 80'h3FFA_FFAADDB967EF5000; // atan(2^- 4) = 0.06241880999595735002 rad ( 3.57633°)
            6'd 5: atan_value = 80'h3FF9_FFEAADDD4BB12800; // atan(2^- 5) = 0.03123983343026827744 rad ( 1.78991°)
            6'd 6: atan_value = 80'h3FF8_FFFAAADDDB94D800; // atan(2^- 6) = 0.01562372862047683129 rad ( 0.89517°)
            6'd 7: atan_value = 80'h3FF7_FFFEAAADDDD4B800; // atan(2^- 7) = 0.00781234106010111114 rad ( 0.44761°)
            6'd 8: atan_value = 80'h3FF6_FFFFAAAADDDDB800; // atan(2^- 8) = 0.00390623013196697176 rad ( 0.22381°)
            6'd 9: atan_value = 80'h3FF5_FFFFEAAAADDDE000; // atan(2^- 9) = 0.00195312251647881876 rad ( 0.11191°)
            6'd10: atan_value = 80'h3FF4_FFFFFAAAAADDE000; // atan(2^-10) = 0.00097656218955931946 rad ( 0.05595°)
            6'd11: atan_value = 80'h3FF3_FFFFFEAAAAADE000; // atan(2^-11) = 0.00048828121119489829 rad ( 0.02798°)
            6'd12: atan_value = 80'h3FF2_FFFFFFAAAAAAE000; // atan(2^-12) = 0.00024414062014936177 rad ( 0.01399°)
            6'd13: atan_value = 80'h3FF1_FFFFFFEAAAAAB000; // atan(2^-13) = 0.00012207031189367021 rad ( 0.00699°)
            6'd14: atan_value = 80'h3FF0_FFFFFFFAAAAAA800; // atan(2^-14) = 0.00006103515617420877 rad ( 0.00350°)
            6'd15: atan_value = 80'h3FEF_FFFFFFFEAAAAA800; // atan(2^-15) = 0.00003051757811552610 rad ( 0.00175°)
            6'd16: atan_value = 80'h3FEE_FFFFFFFFAAAAA800; // atan(2^-16) = 0.00001525878906131576 rad ( 0.00087°)
            6'd17: atan_value = 80'h3FED_FFFFFFFFEAAAA800; // atan(2^-17) = 0.00000762939453110197 rad ( 0.00044°)
            6'd18: atan_value = 80'h3FEC_FFFFFFFFFAAAA800; // atan(2^-18) = 0.00000381469726560650 rad ( 0.00022°)
            6'd19: atan_value = 80'h3FEB_FFFFFFFFFEAAA800; // atan(2^-19) = 0.00000190734863281019 rad ( 0.00011°)
            6'd20: atan_value = 80'h3FEA_FFFFFFFFFFAAA800; // atan(2^-20) = 0.00000095367431640596 rad ( 0.00005°)
            6'd21: atan_value = 80'h3FE9_FFFFFFFFFFEAA800; // atan(2^-21) = 0.00000047683715820309 rad ( 0.00003°)
            6'd22: atan_value = 80'h3FE8_FFFFFFFFFFFAA800; // atan(2^-22) = 0.00000023841857910156 rad ( 0.00001°)
            6'd23: atan_value = 80'h3FE7_FFFFFFFFFFFEA800; // atan(2^-23) = 0.00000011920928955078 rad ( 0.00001°)
            6'd24: atan_value = 80'h3FE7_7FFFFFFFFFFFD400; // atan(2^-24) = 0.00000005960464477539 rad ( 0.00000°)
            6'd25: atan_value = 80'h3FE6_7FFFFFFFFFFFF400; // atan(2^-25) = 0.00000002980232238770 rad ( 0.00000°)
            6'd26: atan_value = 80'h3FE5_7FFFFFFFFFFFFC00; // atan(2^-26) = 0.00000001490116119385 rad ( 0.00000°)
            6'd27: atan_value = 80'h3FE4_8000000000000000; // atan(2^-27) = 0.00000000745058059692 rad ( 0.00000°)
            6'd28: atan_value = 80'h3FE3_8000000000000000; // atan(2^-28) = 0.00000000372529029846 rad ( 0.00000°)
            6'd29: atan_value = 80'h3FE2_8000000000000000; // atan(2^-29) = 0.00000000186264514923 rad ( 0.00000°)
            6'd30: atan_value = 80'h3FE1_8000000000000000; // atan(2^-30) = 0.00000000093132257462 rad ( 0.00000°)
            6'd31: atan_value = 80'h3FE0_8000000000000000; // atan(2^-31) = 0.00000000046566128731 rad ( 0.00000°)
            6'd32: atan_value = 80'h3FDF_8000000000000000; // atan(2^-32) = 0.00000000023283064365 rad ( 0.00000°)
            6'd33: atan_value = 80'h3FDE_8000000000000000; // atan(2^-33) = 0.00000000011641532183 rad ( 0.00000°)
            6'd34: atan_value = 80'h3FDD_8000000000000000; // atan(2^-34) = 0.00000000005820766091 rad ( 0.00000°)
            6'd35: atan_value = 80'h3FDC_8000000000000000; // atan(2^-35) = 0.00000000002910383046 rad ( 0.00000°)
            6'd36: atan_value = 80'h3FDB_8000000000000000; // atan(2^-36) = 0.00000000001455191523 rad ( 0.00000°)
            6'd37: atan_value = 80'h3FDA_8000000000000000; // atan(2^-37) = 0.00000000000727595761 rad ( 0.00000°)
            6'd38: atan_value = 80'h3FD9_8000000000000000; // atan(2^-38) = 0.00000000000363797881 rad ( 0.00000°)
            6'd39: atan_value = 80'h3FD8_8000000000000000; // atan(2^-39) = 0.00000000000181898940 rad ( 0.00000°)
            6'd40: atan_value = 80'h3FD7_8000000000000000; // atan(2^-40) = 0.00000000000090949470 rad ( 0.00000°)
            6'd41: atan_value = 80'h3FD6_8000000000000000; // atan(2^-41) = 0.00000000000045474735 rad ( 0.00000°)
            6'd42: atan_value = 80'h3FD5_8000000000000000; // atan(2^-42) = 0.00000000000022737368 rad ( 0.00000°)
            6'd43: atan_value = 80'h3FD4_8000000000000000; // atan(2^-43) = 0.00000000000011368684 rad ( 0.00000°)
            6'd44: atan_value = 80'h3FD3_8000000000000000; // atan(2^-44) = 0.00000000000005684342 rad ( 0.00000°)
            6'd45: atan_value = 80'h3FD2_8000000000000000; // atan(2^-45) = 0.00000000000002842171 rad ( 0.00000°)
            6'd46: atan_value = 80'h3FD1_8000000000000000; // atan(2^-46) = 0.00000000000001421085 rad ( 0.00000°)
            6'd47: atan_value = 80'h3FD0_8000000000000000; // atan(2^-47) = 0.00000000000000710543 rad ( 0.00000°)
            6'd48: atan_value = 80'h3FCF_8000000000000000; // atan(2^-48) = 0.00000000000000355271 rad ( 0.00000°)
            6'd49: atan_value = 80'h3FCE_8000000000000000; // atan(2^-49) = 0.00000000000000177636 rad ( 0.00000°)
            6'd50: atan_value = 80'h3FCD_8000000000000000; // atan(2^-50) = 0.00000000000000088818 rad ( 0.00000°)
            6'd51: atan_value = 80'h3FCC_8000000000000000; // atan(2^-51) = 0.00000000000000044409 rad ( 0.00000°)
            6'd52: atan_value = 80'h3FCB_8000000000000000; // atan(2^-52) = 0.00000000000000022204 rad ( 0.00000°)
            6'd53: atan_value = 80'h3FCA_8000000000000000; // atan(2^-53) = 0.00000000000000011102 rad ( 0.00000°)
            6'd54: atan_value = 80'h3FC9_8000000000000000; // atan(2^-54) = 0.00000000000000005551 rad ( 0.00000°)
            6'd55: atan_value = 80'h3FC8_8000000000000000; // atan(2^-55) = 0.00000000000000002776 rad ( 0.00000°)
            6'd56: atan_value = 80'h3FC7_8000000000000000; // atan(2^-56) = 0.00000000000000001388 rad ( 0.00000°)
            6'd57: atan_value = 80'h3FC6_8000000000000000; // atan(2^-57) = 0.00000000000000000694 rad ( 0.00000°)
            6'd58: atan_value = 80'h3FC5_8000000000000000; // atan(2^-58) = 0.00000000000000000347 rad ( 0.00000°)
            6'd59: atan_value = 80'h3FC4_8000000000000000; // atan(2^-59) = 0.00000000000000000173 rad ( 0.00000°)
            6'd60: atan_value = 80'h3FC3_8000000000000000; // atan(2^-60) = 0.00000000000000000087 rad ( 0.00000°)
            6'd61: atan_value = 80'h3FC2_8000000000000000; // atan(2^-61) = 0.00000000000000000043 rad ( 0.00000°)
            6'd62: atan_value = 80'h3FC1_8000000000000000; // atan(2^-62) = 0.00000000000000000022 rad ( 0.00000°)
            6'd63: atan_value = 80'h3FC0_8000000000000000; // atan(2^-63) = 0.00000000000000000011 rad ( 0.00000°)
            default: atan_value = 80'h0; // Should never occur
        endcase
    end

endmodule

//=====================================================================
// Verification Notes
//=====================================================================
//
// Key values for reference:
//
// atan(2^- 0) = 0.78539816339744827900 rad
// atan(2^- 1) = 0.46364760900080609352 rad
// atan(2^- 2) = 0.24497866312686414347 rad
// atan(2^- 3) = 0.12435499454676143816 rad
// atan(2^- 4) = 0.06241880999595735002 rad
// atan(2^-10) = 0.00097656218955931946 rad
// atan(2^-20) = 0.00000095367431640596 rad
// atan(2^-30) = 0.00000000093132257462 rad
// atan(2^-40) = 0.00000000000090949470 rad
// atan(2^-50) = 0.00000000000000088818 rad
// atan(2^-63) = 0.00000000000000000011 rad
//
// The convergence domain of CORDIC is approximately [-99.7°, +99.7°]
// or [-1.74 rad, +1.74 rad].
//
// For angles outside this range, use range reduction:
// - Map to [-π, π] using modulo 2π
// - Use trig identities to map to [-π/4, π/4] for best accuracy
//
// Sum of all atan values ≈ 1.74328 radians ≈ 99.88°
// This represents the maximum angle that can be reduced to zero
// in rotation mode CORDIC.
//=====================================================================
