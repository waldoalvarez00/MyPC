// Copyright 2025, Waldo Alvarez, https://pipflow.com
//
// Comprehensive Testbench for Pipelined Arbiters
// Tests PipelinedDMAArbiter and PipelinedMemArbiterExtend
// Fixed memory model timing for proper pipelined operation
//
//============================================================================

`timescale 1ns/1ps
`default_nettype none

module pipelined_arbiters_comprehensive_tb;

//============================================================================
// Test Configuration
//============================================================================

parameter CLK_PERIOD = 20;  // 50 MHz
parameter MEM_LATENCY = 3;  // SDRAM latency in cycles

//============================================================================
// Test 1: PipelinedDMAArbiter
//============================================================================

reg clk, reset;

// DMA bus (A-bus)
reg  [19:1] dma_addr;
wire [15:0] dma_data_in;
reg  [15:0] dma_data_out;
reg         dma_access;
wire        dma_ack;
reg         dma_wr_en;
reg  [1:0]  dma_bytesel;

// CPU bus (B-bus)
reg  [19:1] cpu_addr;
wire [15:0] cpu_data_in;
reg  [15:0] cpu_data_out;
reg         cpu_access;
wire        cpu_ack;
reg         cpu_wr_en;
reg  [1:0]  cpu_bytesel;

// Memory interface from DMA arbiter
wire [19:1] mem_addr_dma;
reg  [15:0] mem_data_in_dma;
wire [15:0] mem_data_out_dma;
wire        mem_access_dma;
reg         mem_ack_dma;
wire        mem_wr_en_dma;
wire [1:0]  mem_bytesel_dma;

// Test tracking
integer test_num;
integer pass_count;
integer fail_count;
integer cycle_count;

// Memory model
reg [15:0] memory [0:524287];

// DUT 1: PipelinedDMAArbiter
PipelinedDMAArbiter dma_arbiter (
    .clk(clk),
    .reset(reset),
    // A-bus (DMA)
    .a_m_addr(dma_addr),
    .a_m_data_in(dma_data_in),
    .a_m_data_out(dma_data_out),
    .a_m_access(dma_access),
    .a_m_ack(dma_ack),
    .a_m_wr_en(dma_wr_en),
    .a_m_bytesel(dma_bytesel),
    .ioa(1'b0),
    // B-bus (CPU)
    .b_m_addr(cpu_addr),
    .b_m_data_in(cpu_data_in),
    .b_m_data_out(cpu_data_out),
    .b_m_access(cpu_access),
    .b_m_ack(cpu_ack),
    .b_m_wr_en(cpu_wr_en),
    .b_m_bytesel(cpu_bytesel),
    .iob(1'b0),
    // Output
    .q_m_addr(mem_addr_dma),
    .q_m_data_in(mem_data_in_dma),
    .q_m_data_out(mem_data_out_dma),
    .q_m_access(mem_access_dma),
    .q_m_ack(mem_ack_dma),
    .q_m_wr_en(mem_wr_en_dma),
    .q_m_bytesel(mem_bytesel_dma),
    .ioq(),
    .q_b()
);

//============================================================================
// Test 2: PipelinedMemArbiterExtend
//============================================================================

// CPU+DMA bus
reg  [19:1] cpudma_addr;
wire [15:0] cpudma_data_in;
reg  [15:0] cpudma_data_out;
reg         cpudma_access;
wire        cpudma_ack;
reg         cpudma_wr_en;
reg  [1:0]  cpudma_bytesel;

// VGA bus
reg  [19:1] vga_addr;
wire [15:0] vga_data_in;
reg  [15:0] vga_data_out;
reg         vga_access;
wire        vga_ack;
reg         vga_wr_en;
reg  [1:0]  vga_bytesel;

// VGA priority
reg vga_active_display;

// SDRAM interface from mem arbiter
wire [19:1] sdram_addr;
reg  [15:0] sdram_data_in;
wire [15:0] sdram_data_out;
wire        sdram_access;
reg         sdram_ack;
wire        sdram_wr_en;
wire [1:0]  sdram_bytesel;

// DUT 2: PipelinedMemArbiterExtend
PipelinedMemArbiterExtend mem_arbiter (
    .clk(clk),
    .reset(reset),
    // CPU+DMA bus
    .cpu_m_addr(cpudma_addr),
    .cpu_m_data_in(cpudma_data_in),
    .cpu_m_data_out(cpudma_data_out),
    .cpu_m_access(cpudma_access),
    .cpu_m_ack(cpudma_ack),
    .cpu_m_wr_en(cpudma_wr_en),
    .cpu_m_bytesel(cpudma_bytesel),
    // VGA bus
    .mcga_m_addr(vga_addr),
    .mcga_m_data_in(vga_data_in),
    .mcga_m_data_out(vga_data_out),
    .mcga_m_access(vga_access),
    .mcga_m_ack(vga_ack),
    .mcga_m_wr_en(vga_wr_en),
    .mcga_m_bytesel(vga_bytesel),
    // Priority hint
    .vga_active_display(vga_active_display),
    // SDRAM
    .sdram_m_addr(sdram_addr),
    .sdram_m_data_in(sdram_data_in),
    .sdram_m_data_out(sdram_data_out),
    .sdram_m_access(sdram_access),
    .sdram_m_ack(sdram_ack),
    .sdram_m_wr_en(sdram_wr_en),
    .sdram_m_bytesel(sdram_bytesel),
    .q_b()
);

//============================================================================
// Clock Generation
//============================================================================

initial begin
    clk = 0;
    forever #(CLK_PERIOD/2) clk = ~clk;
end

//============================================================================
// Memory Model - Improved Timing for Pipelined Operation
//============================================================================

// Memory model for DMA arbiter output
integer mem_dma_latency_counter;
reg mem_dma_pending;

always @(posedge clk) begin
    if (reset) begin
        mem_ack_dma <= 1'b0;
        mem_dma_latency_counter <= 0;
        mem_dma_pending <= 1'b0;
    end else begin
        if (mem_access_dma && !mem_dma_pending) begin
            // New request
            mem_dma_pending <= 1'b1;
            mem_dma_latency_counter <= MEM_LATENCY;
            mem_ack_dma <= 1'b0;
        end else if (mem_dma_pending) begin
            if (mem_dma_latency_counter > 1) begin
                mem_dma_latency_counter <= mem_dma_latency_counter - 1;
                mem_ack_dma <= 1'b0;
            end else begin
                // Acknowledge
                mem_ack_dma <= 1'b1;
                mem_dma_pending <= 1'b0;
                // Handle read/write
                if (mem_wr_en_dma) begin
                    memory[mem_addr_dma] <= mem_data_out_dma;
                end else begin
                    mem_data_in_dma <= memory[mem_addr_dma];
                end
            end
        end else begin
            mem_ack_dma <= 1'b0;
        end
    end
end

// Memory model for mem arbiter output
integer sdram_latency_counter;
reg sdram_pending;

always @(posedge clk) begin
    if (reset) begin
        sdram_ack <= 1'b0;
        sdram_latency_counter <= 0;
        sdram_pending <= 1'b0;
    end else begin
        if (sdram_access && !sdram_pending) begin
            // New request
            sdram_pending <= 1'b1;
            sdram_latency_counter <= MEM_LATENCY;
            sdram_ack <= 1'b0;
        end else if (sdram_pending) begin
            if (sdram_latency_counter > 1) begin
                sdram_latency_counter <= sdram_latency_counter - 1;
                sdram_ack <= 1'b0;
            end else begin
                // Acknowledge
                sdram_ack <= 1'b1;
                sdram_pending <= 1'b0;
                // Handle read/write
                if (sdram_wr_en) begin
                    memory[sdram_addr] <= sdram_data_out;
                end else begin
                    sdram_data_in <= memory[sdram_addr];
                end
            end
        end else begin
            sdram_ack <= 1'b0;
        end
    end
end

//============================================================================
// Test Utilities
//============================================================================

task check_result(input condition, input string description);
begin
    test_num = test_num + 1;
    if (condition) begin
        pass_count = pass_count + 1;
        $display("  [PASS] Test %0d: %s", test_num, description);
    end else begin
        fail_count = fail_count + 1;
        $display("  [FAIL] Test %0d: %s", test_num, description);
    end
end
endtask

task init_memory();
    integer i;
begin
    for (i = 0; i < 524288; i = i + 1) begin
        memory[i] = i[15:0] ^ 16'hA5A5;
    end
end
endtask

//============================================================================
// Main Test Sequence
//============================================================================

initial begin
    // Initialize
    test_num = 0;
    pass_count = 0;
    fail_count = 0;
    cycle_count = 0;

    reset = 1;
    dma_access = 0;
    cpu_access = 0;
    cpudma_access = 0;
    vga_access = 0;
    dma_wr_en = 0;
    cpu_wr_en = 0;
    cpudma_wr_en = 0;
    vga_wr_en = 0;
    vga_active_display = 0;

    $display("========================================");
    $display("Comprehensive Pipelined Arbiters Test");
    $display("========================================\n");

    init_memory();

    repeat(10) @(posedge clk);
    reset = 0;
    repeat(5) @(posedge clk);

    //========================================================================
    // TEST SUITE 1: PipelinedDMAArbiter
    //========================================================================

    $display("TEST SUITE 1: PipelinedDMAArbiter");
    $display("----------------------------------\n");

    // Test 1.1: Basic CPU read
    $display("Test 1.1: Basic CPU read");
    cpu_addr = 19'h01000;
    cpu_data_out = 16'h0000;
    cpu_wr_en = 1'b0;
    cpu_bytesel = 2'b11;
    cpu_access = 1'b1;

    @(posedge clk);
    wait(cpu_ack);
    check_result(cpu_data_in == (16'h1000 ^ 16'hA5A5), "CPU read data correct");
    cpu_access = 1'b0;
    @(posedge clk);

    // Test 1.2: Basic DMA read
    $display("\nTest 1.2: Basic DMA read");
    dma_addr = 19'h02000;
    dma_data_out = 16'h0000;
    dma_wr_en = 1'b0;
    dma_bytesel = 2'b11;
    dma_access = 1'b1;

    @(posedge clk);
    wait(dma_ack);
    check_result(dma_data_in == (16'h2000 ^ 16'hA5A5), "DMA read data correct");
    dma_access = 1'b0;
    @(posedge clk);

    // Test 1.3: CPU priority (both request)
    $display("\nTest 1.3: CPU priority when both request");
    fork
        begin
            dma_addr = 19'h03000;
            dma_access = 1'b1;
            dma_wr_en = 1'b0;
            dma_bytesel = 2'b11;
        end
        begin
            cpu_addr = 19'h04000;
            cpu_access = 1'b1;
            cpu_wr_en = 1'b0;
            cpu_bytesel = 2'b11;
        end
    join

    @(posedge clk);
    wait(cpu_ack || dma_ack);
    check_result(cpu_ack && !dma_ack, "CPU has priority");
    wait(dma_ack);
    check_result(dma_ack, "DMA served after CPU");
    dma_access = 1'b0;
    cpu_access = 1'b0;
    @(posedge clk);

    // Test 1.4: Write operations
    $display("\nTest 1.4: Write operations");
    cpu_addr = 19'h05000;
    cpu_data_out = 16'hDEAD;
    cpu_wr_en = 1'b1;
    cpu_bytesel = 2'b11;
    cpu_access = 1'b1;

    @(posedge clk);
    wait(cpu_ack);
    cpu_access = 1'b0;
    cpu_wr_en = 1'b0;
    @(posedge clk);

    // Read back
    cpu_addr = 19'h05000;
    cpu_wr_en = 1'b0;
    cpu_access = 1'b1;
    @(posedge clk);
    wait(cpu_ack);
    check_result(cpu_data_in == 16'hDEAD, "CPU write verified");
    cpu_access = 1'b0;
    @(posedge clk);

    // Test 1.5: Back-to-back throughput
    $display("\nTest 1.5: Back-to-back throughput test");
    begin
        integer start_cycle, end_cycle, i;
        real throughput;

        start_cycle = cycle_count;

        for (i = 0; i < 20; i = i + 1) begin
            cpu_addr = 19'h10000 + i;
            cpu_wr_en = 1'b0;
            cpu_bytesel = 2'b11;
            cpu_access = 1'b1;
            @(posedge clk);
            wait(cpu_ack);
            cpu_access = 1'b0;
            @(posedge clk);
        end

        end_cycle = cycle_count;
        throughput = real'(20) / real'(end_cycle - start_cycle);

        $display("  20 operations in %0d cycles", end_cycle - start_cycle);
        $display("  Throughput: %.3f ops/cycle", throughput);
        check_result(throughput >= 0.30,
                    $sformatf("Throughput %.3f >= 0.30", throughput));
    end

    //========================================================================
    // TEST SUITE 2: PipelinedMemArbiterExtend
    //========================================================================

    $display("\n\nTEST SUITE 2: PipelinedMemArbiterExtend");
    $display("----------------------------------------\n");

    // Test 2.1: Basic CPU+DMA read
    $display("Test 2.1: Basic CPU+DMA read");
    cpudma_addr = 19'h01000;
    cpudma_data_out = 16'h0000;
    cpudma_wr_en = 1'b0;
    cpudma_bytesel = 2'b11;
    cpudma_access = 1'b1;

    @(posedge clk);
    wait(cpudma_ack);
    check_result(cpudma_data_in == (16'h1000 ^ 16'hA5A5), "CPU+DMA read data correct");
    cpudma_access = 1'b0;
    @(posedge clk);

    // Test 2.2: Basic VGA read
    $display("\nTest 2.2: Basic VGA read");
    vga_addr = 19'h02000;
    vga_data_out = 16'h0000;
    vga_wr_en = 1'b0;
    vga_bytesel = 2'b11;
    vga_access = 1'b1;

    @(posedge clk);
    wait(vga_ack);
    check_result(vga_data_in == (16'h2000 ^ 16'hA5A5), "VGA read data correct");
    vga_access = 1'b0;
    @(posedge clk);

    // Test 2.3: VGA priority during active display
    $display("\nTest 2.3: VGA priority during active display");
    vga_active_display = 1'b1;

    fork
        begin
            cpudma_addr = 19'h03000;
            cpudma_access = 1'b1;
            cpudma_wr_en = 1'b0;
            cpudma_bytesel = 2'b11;
        end
        begin
            vga_addr = 19'h04000;
            vga_access = 1'b1;
            vga_wr_en = 1'b0;
            vga_bytesel = 2'b11;
        end
    join

    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    wait(vga_ack || cpudma_ack);
    check_result(vga_ack && !cpudma_ack, "VGA has priority during active display");
    wait(cpudma_ack);
    check_result(cpudma_ack, "CPU+DMA served after VGA");
    cpudma_access = 1'b0;
    vga_access = 1'b0;
    vga_active_display = 1'b0;
    @(posedge clk);

    // Test 2.4: Write operations
    $display("\nTest 2.4: Write operations");
    cpudma_addr = 19'h05000;
    cpudma_data_out = 16'hBEEF;
    cpudma_wr_en = 1'b1;
    cpudma_bytesel = 2'b11;
    cpudma_access = 1'b1;

    @(posedge clk);
    wait(cpudma_ack);
    cpudma_access = 1'b0;
    cpudma_wr_en = 1'b0;
    @(posedge clk);

    // Read back
    cpudma_addr = 19'h05000;
    cpudma_wr_en = 1'b0;
    cpudma_access = 1'b1;
    @(posedge clk);
    wait(cpudma_ack);
    check_result(cpudma_data_in == 16'hBEEF, "CPU+DMA write verified");
    cpudma_access = 1'b0;
    @(posedge clk);

    // Test 2.5: Interleaved requests
    $display("\nTest 2.5: Interleaved CPU+DMA and VGA requests");
    begin
        integer i;

        for (i = 0; i < 10; i = i + 1) begin
            // CPU+DMA request
            cpudma_addr = 19'h10000 + i;
            cpudma_wr_en = 1'b0;
            cpudma_bytesel = 2'b11;
            cpudma_access = 1'b1;
            @(posedge clk);
            wait(cpudma_ack);
            cpudma_access = 1'b0;
            @(posedge clk);

            // VGA request
            vga_addr = 19'h20000 + i;
            vga_wr_en = 1'b0;
            vga_bytesel = 2'b11;
            vga_access = 1'b1;
            @(posedge clk);
            wait(vga_ack);
            vga_access = 1'b0;
            @(posedge clk);
        end

        check_result(1, "Interleaved requests completed");
    end

    // Test 2.6: Fairness test
    $display("\nTest 2.6: Round-robin fairness test");
    begin
        integer vga_first, cpu_first, i;
        vga_first = 0;
        cpu_first = 0;

        vga_active_display = 1'b0;  // No priority

        for (i = 0; i < 10; i = i + 1) begin
            fork
                begin
                    cpudma_addr = 19'h30000 + i;
                    cpudma_access = 1'b1;
                    cpudma_wr_en = 1'b0;
                    cpudma_bytesel = 2'b11;
                end
                begin
                    vga_addr = 19'h40000 + i;
                    vga_access = 1'b1;
                    vga_wr_en = 1'b0;
                    vga_bytesel = 2'b11;
                end
            join

            @(posedge clk);
            @(posedge clk);
            @(posedge clk);
            @(posedge clk);

            if (cpudma_ack) cpu_first = cpu_first + 1;
            if (vga_ack) vga_first = vga_first + 1;

            wait(cpudma_ack && vga_ack);
            cpudma_access = 1'b0;
            vga_access = 1'b0;
            @(posedge clk);
        end

        $display("  CPU+DMA served first: %0d times", cpu_first);
        $display("  VGA served first: %0d times", vga_first);
        check_result(cpu_first >= 3 && vga_first >= 3, "Fair round-robin arbitration");
    end

    //========================================================================
    // Test Summary
    //========================================================================

    repeat(10) @(posedge clk);

    $display("\n========================================");
    $display("TEST SUMMARY");
    $display("========================================");
    $display("Total tests: %0d", test_num);
    $display("Passed:      %0d", pass_count);
    $display("Failed:      %0d", fail_count);
    $display("Success rate: %.1f%%", real'(pass_count) / real'(test_num) * 100.0);
    $display("========================================\n");

    if (fail_count == 0) begin
        $display("*** ALL TESTS PASSED ***\n");
        $finish(0);
    end else begin
        $display("*** SOME TESTS FAILED ***\n");
        $finish(1);
    end
end

// Cycle counter
always @(posedge clk) begin
    if (!reset) cycle_count <= cycle_count + 1;
end

// Timeout watchdog
initial begin
    #1000000;  // 1ms timeout
    $display("\n========================================");
    $display("ERROR: Simulation timeout!");
    $display("========================================");
    $finish(2);
end

// Waveform dump
initial begin
    $dumpfile("pipelined_arbiters_comprehensive_tb.vcd");
    $dumpvars(0, pipelined_arbiters_comprehensive_tb);
end

endmodule
`default_nettype wire
