// Copyright Jamie Iles, 2018
//
// This file is part of s80x86.
//
// s80x86 is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// s80x86 is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with s80x86.  If not, see <http://www.gnu.org/licenses/>.

function logic insn_has_modrm;
    input logic [7:0] opcode;

    casez (opcode)
    8'h87: insn_has_modrm = 1'b1;
    8'h8a: insn_has_modrm = 1'b1;
    8'hd2: insn_has_modrm = 1'b1;
    8'h21: insn_has_modrm = 1'b1;
    8'h86: insn_has_modrm = 1'b1;
    8'h19: insn_has_modrm = 1'b1;
    8'hdb: insn_has_modrm = 1'b1;
    8'h84: insn_has_modrm = 1'b1;
    8'hdf: insn_has_modrm = 1'b1;
    8'hd1: insn_has_modrm = 1'b1;
    8'h31: insn_has_modrm = 1'b1;
    8'h89: insn_has_modrm = 1'b1;
    8'h28: insn_has_modrm = 1'b1;
    8'h62: insn_has_modrm = 1'b1;
    8'hd0: insn_has_modrm = 1'b1;
    8'h29: insn_has_modrm = 1'b1;
    8'h2a: insn_has_modrm = 1'b1;
    8'h09: insn_has_modrm = 1'b1;
    8'hd3: insn_has_modrm = 1'b1;
    8'h22: insn_has_modrm = 1'b1;
    8'hd9: insn_has_modrm = 1'b1;
    8'h1b: insn_has_modrm = 1'b1;
    8'h33: insn_has_modrm = 1'b1;
    8'h12: insn_has_modrm = 1'b1;
    8'h1a: insn_has_modrm = 1'b1;
    8'hdd: insn_has_modrm = 1'b1;
    8'hdc: insn_has_modrm = 1'b1;
    8'h6b: insn_has_modrm = 1'b1;
    8'hf6: insn_has_modrm = 1'b1;
    8'h30: insn_has_modrm = 1'b1;
    8'h13: insn_has_modrm = 1'b1;
    8'hfe: insn_has_modrm = 1'b1;
    8'h8e: insn_has_modrm = 1'b1;
    8'h85: insn_has_modrm = 1'b1;
    8'h39: insn_has_modrm = 1'b1;
    8'h20: insn_has_modrm = 1'b1;
    8'h23: insn_has_modrm = 1'b1;
    8'hf7: insn_has_modrm = 1'b1;
    8'h10: insn_has_modrm = 1'b1;
    8'h0a: insn_has_modrm = 1'b1;
    8'h01: insn_has_modrm = 1'b1;
    8'h08: insn_has_modrm = 1'b1;
    8'h81: insn_has_modrm = 1'b1;
    8'h11: insn_has_modrm = 1'b1;
    8'hc7: insn_has_modrm = 1'b1;
    8'h32: insn_has_modrm = 1'b1;
    8'h8d: insn_has_modrm = 1'b1;
    8'h83: insn_has_modrm = 1'b1;
    8'h03: insn_has_modrm = 1'b1;
    8'h8b: insn_has_modrm = 1'b1;
    8'h0b: insn_has_modrm = 1'b1;
    8'hc6: insn_has_modrm = 1'b1;
    8'h3a: insn_has_modrm = 1'b1;
    8'h18: insn_has_modrm = 1'b1;
    8'h80: insn_has_modrm = 1'b1;
    8'hc5: insn_has_modrm = 1'b1;
    8'h00: insn_has_modrm = 1'b1;
    8'h3b: insn_has_modrm = 1'b1;
    8'hc0: insn_has_modrm = 1'b1;
    8'hde: insn_has_modrm = 1'b1;
    8'hd8: insn_has_modrm = 1'b1;
    8'h69: insn_has_modrm = 1'b1;
    8'h8c: insn_has_modrm = 1'b1;
    8'h2b: insn_has_modrm = 1'b1;
    8'h02: insn_has_modrm = 1'b1;
    8'hff: insn_has_modrm = 1'b1;
    8'h88: insn_has_modrm = 1'b1;
    8'hda: insn_has_modrm = 1'b1;
    8'h82: insn_has_modrm = 1'b1;
    8'hc4: insn_has_modrm = 1'b1;
    8'h38: insn_has_modrm = 1'b1;
    8'h8f: insn_has_modrm = 1'b1;
    8'hc1: insn_has_modrm = 1'b1;
    default: insn_has_modrm = 1'b0;
    endcase
endfunction

function logic [1:0] insn_immed_count;
    input logic [7:0] opcode;
    input logic [2:0] modrm_reg;

    unique casez ({opcode, modrm_reg})
    {8'h37, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hd5, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hd4, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h3f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h10, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h11, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h12, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h13, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h14, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h15, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h2}: insn_immed_count = 2'd1;
    {8'h81, 3'h2}: insn_immed_count = 2'd1;
    {8'h82, 3'h2}: insn_immed_count = 2'd1;
    {8'h83, 3'h2}: insn_immed_count = 2'd1;
    {8'h00, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h01, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h02, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h03, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h04, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h05, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h0}: insn_immed_count = 2'd1;
    {8'h81, 3'h0}: insn_immed_count = 2'd1;
    {8'h82, 3'h0}: insn_immed_count = 2'd1;
    {8'h83, 3'h0}: insn_immed_count = 2'd1;
    {8'h20, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h21, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h22, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h23, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h24, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h25, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h4}: insn_immed_count = 2'd1;
    {8'h81, 3'h4}: insn_immed_count = 2'd1;
    {8'h82, 3'h4}: insn_immed_count = 2'd1;
    {8'h83, 3'h4}: insn_immed_count = 2'd1;
    {8'h62, 3'bzzz}: insn_immed_count = 2'd0;
    {8'he8, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h9a, 3'bzzz}: insn_immed_count = 2'd2;
    {8'hff, 3'h2}: insn_immed_count = 2'd0;
    {8'hff, 3'h3}: insn_immed_count = 2'd0;
    {8'h98, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hf8, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hfc, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hfa, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hf5, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h38, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h39, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h3a, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h3b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h3c, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h3d, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h7}: insn_immed_count = 2'd1;
    {8'h81, 3'h7}: insn_immed_count = 2'd1;
    {8'h82, 3'h7}: insn_immed_count = 2'd1;
    {8'h83, 3'h7}: insn_immed_count = 2'd1;
    {8'ha6, 3'bzzz}: insn_immed_count = 2'd0;
    {8'ha7, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h99, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h27, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h2f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hfe, 3'h1}: insn_immed_count = 2'd0;
    {8'hff, 3'h1}: insn_immed_count = 2'd0;
    {8'h48, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h49, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h4a, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h4b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h4c, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h4d, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h4e, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h4f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hf6, 3'h6}: insn_immed_count = 2'd0;
    {8'hf7, 3'h6}: insn_immed_count = 2'd0;
    {8'hc8, 3'bzzz}: insn_immed_count = 2'd2;
    {8'hd8, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hd9, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hda, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hdb, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hdc, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hdd, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hde, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hdf, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hf4, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hf6, 3'h7}: insn_immed_count = 2'd0;
    {8'hf7, 3'h7}: insn_immed_count = 2'd0;
    {8'hf6, 3'h5}: insn_immed_count = 2'd0;
    {8'hf7, 3'h5}: insn_immed_count = 2'd0;
    {8'h69, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h6b, 3'bzzz}: insn_immed_count = 2'd1;
    {8'he4, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hec, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hfe, 3'h0}: insn_immed_count = 2'd0;
    {8'hff, 3'h0}: insn_immed_count = 2'd0;
    {8'h40, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h41, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h42, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h43, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h44, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h45, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h46, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h47, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h6c, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h6d, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hcd, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hcc, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hce, 3'bzzz}: insn_immed_count = 2'd0;
    {8'he5, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hed, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hcf, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h72, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h76, 3'bzzz}: insn_immed_count = 2'd1;
    {8'he3, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h74, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h7c, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h7e, 3'bzzz}: insn_immed_count = 2'd1;
    {8'he9, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hea, 3'bzzz}: insn_immed_count = 2'd2;
    {8'heb, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hff, 3'h4}: insn_immed_count = 2'd0;
    {8'hff, 3'h5}: insn_immed_count = 2'd0;
    {8'h73, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h77, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h75, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h7d, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h7f, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h71, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h7b, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h79, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h70, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h7a, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h78, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h9f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hc5, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h8d, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hc9, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hc4, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hac, 3'bzzz}: insn_immed_count = 2'd0;
    {8'had, 3'bzzz}: insn_immed_count = 2'd0;
    {8'he2, 3'bzzz}: insn_immed_count = 2'd1;
    {8'he1, 3'bzzz}: insn_immed_count = 2'd1;
    {8'he0, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h88, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h89, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h8a, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h8b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hc6, 3'h0}: insn_immed_count = 2'd1;
    {8'hc7, 3'h0}: insn_immed_count = 2'd1;
    {8'hb0, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb1, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb2, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb3, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb4, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb5, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb6, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb7, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb8, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hb9, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hba, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hbb, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hbc, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hbd, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hbe, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hbf, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h8e, 3'h0}: insn_immed_count = 2'd0;
    {8'h8e, 3'h1}: insn_immed_count = 2'd0;
    {8'h8e, 3'h2}: insn_immed_count = 2'd0;
    {8'h8e, 3'h3}: insn_immed_count = 2'd0;
    {8'h8e, 3'h4}: insn_immed_count = 2'd0;
    {8'h8e, 3'h5}: insn_immed_count = 2'd0;
    {8'h8e, 3'h6}: insn_immed_count = 2'd0;
    {8'h8e, 3'h7}: insn_immed_count = 2'd0;
    {8'h8c, 3'h0}: insn_immed_count = 2'd0;
    {8'h8c, 3'h1}: insn_immed_count = 2'd0;
    {8'h8c, 3'h2}: insn_immed_count = 2'd0;
    {8'h8c, 3'h3}: insn_immed_count = 2'd0;
    {8'h8c, 3'h4}: insn_immed_count = 2'd0;
    {8'h8c, 3'h5}: insn_immed_count = 2'd0;
    {8'h8c, 3'h6}: insn_immed_count = 2'd0;
    {8'h8c, 3'h7}: insn_immed_count = 2'd0;
    {8'ha0, 3'bzzz}: insn_immed_count = 2'd1;
    {8'ha1, 3'bzzz}: insn_immed_count = 2'd1;
    {8'ha2, 3'bzzz}: insn_immed_count = 2'd1;
    {8'ha3, 3'bzzz}: insn_immed_count = 2'd1;
    {8'ha4, 3'bzzz}: insn_immed_count = 2'd0;
    {8'ha5, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hf6, 3'h4}: insn_immed_count = 2'd0;
    {8'hf7, 3'h4}: insn_immed_count = 2'd0;
    {8'hf6, 3'h3}: insn_immed_count = 2'd0;
    {8'hf7, 3'h3}: insn_immed_count = 2'd0;
    {8'h90, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hf6, 3'h2}: insn_immed_count = 2'd0;
    {8'hf7, 3'h2}: insn_immed_count = 2'd0;
    {8'h08, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h09, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h0a, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h0b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h0c, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h0d, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h1}: insn_immed_count = 2'd1;
    {8'h81, 3'h1}: insn_immed_count = 2'd1;
    {8'h82, 3'h1}: insn_immed_count = 2'd1;
    {8'h83, 3'h1}: insn_immed_count = 2'd1;
    {8'he6, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hee, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h6e, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h6f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'he7, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hef, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h58, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h59, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h5a, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h5b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h5c, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h5d, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h5e, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h5f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h07, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h17, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h1f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h8f, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h61, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h9d, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hff, 3'h6}: insn_immed_count = 2'd0;
    {8'h06, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h0e, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h16, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h1e, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h50, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h51, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h52, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h53, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h54, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h55, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h56, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h57, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h68, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h6a, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h60, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h9c, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hd0, 3'h2}: insn_immed_count = 2'd0;
    {8'hd1, 3'h2}: insn_immed_count = 2'd0;
    {8'hc0, 3'h2}: insn_immed_count = 2'd1;
    {8'hc1, 3'h2}: insn_immed_count = 2'd1;
    {8'hd2, 3'h2}: insn_immed_count = 2'd0;
    {8'hd3, 3'h2}: insn_immed_count = 2'd0;
    {8'hd0, 3'h3}: insn_immed_count = 2'd0;
    {8'hd1, 3'h3}: insn_immed_count = 2'd0;
    {8'hc0, 3'h3}: insn_immed_count = 2'd1;
    {8'hc1, 3'h3}: insn_immed_count = 2'd1;
    {8'hd2, 3'h3}: insn_immed_count = 2'd0;
    {8'hd3, 3'h3}: insn_immed_count = 2'd0;
    {8'hc3, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hc2, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hcb, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hca, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hd0, 3'h0}: insn_immed_count = 2'd0;
    {8'hd1, 3'h0}: insn_immed_count = 2'd0;
    {8'hc0, 3'h0}: insn_immed_count = 2'd1;
    {8'hc1, 3'h0}: insn_immed_count = 2'd1;
    {8'hd2, 3'h0}: insn_immed_count = 2'd0;
    {8'hd3, 3'h0}: insn_immed_count = 2'd0;
    {8'hd0, 3'h1}: insn_immed_count = 2'd0;
    {8'hd1, 3'h1}: insn_immed_count = 2'd0;
    {8'hc0, 3'h1}: insn_immed_count = 2'd1;
    {8'hc1, 3'h1}: insn_immed_count = 2'd1;
    {8'hd2, 3'h1}: insn_immed_count = 2'd0;
    {8'hd3, 3'h1}: insn_immed_count = 2'd0;
    {8'h9e, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hd0, 3'h6}: insn_immed_count = 2'd0;
    {8'hd1, 3'h6}: insn_immed_count = 2'd0;
    {8'hc0, 3'h6}: insn_immed_count = 2'd1;
    {8'hc1, 3'h6}: insn_immed_count = 2'd1;
    {8'hd2, 3'h6}: insn_immed_count = 2'd0;
    {8'hd3, 3'h6}: insn_immed_count = 2'd0;
    {8'hd0, 3'h7}: insn_immed_count = 2'd0;
    {8'hd1, 3'h7}: insn_immed_count = 2'd0;
    {8'hc0, 3'h7}: insn_immed_count = 2'd1;
    {8'hc1, 3'h7}: insn_immed_count = 2'd1;
    {8'hd2, 3'h7}: insn_immed_count = 2'd0;
    {8'hd3, 3'h7}: insn_immed_count = 2'd0;
    {8'h18, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h19, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h1a, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h1b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h1c, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h1d, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h3}: insn_immed_count = 2'd1;
    {8'h81, 3'h3}: insn_immed_count = 2'd1;
    {8'h82, 3'h3}: insn_immed_count = 2'd1;
    {8'h83, 3'h3}: insn_immed_count = 2'd1;
    {8'hae, 3'bzzz}: insn_immed_count = 2'd0;
    {8'haf, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hd6, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hd0, 3'h4}: insn_immed_count = 2'd0;
    {8'hd1, 3'h4}: insn_immed_count = 2'd0;
    {8'hc0, 3'h4}: insn_immed_count = 2'd1;
    {8'hc1, 3'h4}: insn_immed_count = 2'd1;
    {8'hd2, 3'h4}: insn_immed_count = 2'd0;
    {8'hd3, 3'h4}: insn_immed_count = 2'd0;
    {8'hd0, 3'h5}: insn_immed_count = 2'd0;
    {8'hd1, 3'h5}: insn_immed_count = 2'd0;
    {8'hc0, 3'h5}: insn_immed_count = 2'd1;
    {8'hc1, 3'h5}: insn_immed_count = 2'd1;
    {8'hd2, 3'h5}: insn_immed_count = 2'd0;
    {8'hd3, 3'h5}: insn_immed_count = 2'd0;
    {8'hf9, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hfd, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hfb, 3'bzzz}: insn_immed_count = 2'd0;
    {8'haa, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hab, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h28, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h29, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h2a, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h2b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h2c, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h2d, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h5}: insn_immed_count = 2'd1;
    {8'h81, 3'h5}: insn_immed_count = 2'd1;
    {8'h82, 3'h5}: insn_immed_count = 2'd1;
    {8'h83, 3'h5}: insn_immed_count = 2'd1;
    {8'h84, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h85, 3'bzzz}: insn_immed_count = 2'd0;
    {8'ha8, 3'bzzz}: insn_immed_count = 2'd1;
    {8'ha9, 3'bzzz}: insn_immed_count = 2'd1;
    {8'hf6, 3'h0}: insn_immed_count = 2'd1;
    {8'hf6, 3'h1}: insn_immed_count = 2'd1;
    {8'hf7, 3'h0}: insn_immed_count = 2'd1;
    {8'hf7, 3'h1}: insn_immed_count = 2'd1;
    {8'h9b, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h86, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h87, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h91, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h92, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h93, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h94, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h95, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h96, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h97, 3'bzzz}: insn_immed_count = 2'd0;
    {8'hd7, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h30, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h31, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h32, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h33, 3'bzzz}: insn_immed_count = 2'd0;
    {8'h34, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h35, 3'bzzz}: insn_immed_count = 2'd1;
    {8'h80, 3'h6}: insn_immed_count = 2'd1;
    {8'h81, 3'h6}: insn_immed_count = 2'd1;
    {8'h82, 3'h6}: insn_immed_count = 2'd1;
    {8'h83, 3'h6}: insn_immed_count = 2'd1;
    default: insn_immed_count = 2'b0;
    endcase
endfunction

function logic insn_immed_is_8bit;
    input logic [7:0] opcode;
    input logic [2:0] modrm_reg;
    input logic immed_num;

    unique casez ({opcode, modrm_reg})
    {8'h37, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd5, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd4, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h3f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h10, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h11, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h12, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h13, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h14, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h15, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h2}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h00, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h01, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h02, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h03, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h04, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h05, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h0}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h20, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h21, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h22, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h23, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h24, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h25, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h4}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h62, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he8, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h9a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h3 & (2'b1 << immed_num));
    {8'hff, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hff, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h98, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf8, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hfc, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hfa, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf5, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h38, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h39, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h3a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h3b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h3c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h3d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h7}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'ha6, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'ha7, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h99, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h27, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h2f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hfe, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hff, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h48, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h49, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h4a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h4b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h4c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h4d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h4e, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h4f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf6, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf7, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc8, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hd8, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd9, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hda, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hdb, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hdc, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hdd, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hde, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hdf, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf4, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf6, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf7, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf6, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf7, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h69, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h6b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he4, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hec, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hfe, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hff, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h40, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h41, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h42, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h43, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h44, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h45, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h46, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h47, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h6c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h6d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hcd, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hcc, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hce, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he5, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hed, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hcf, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h72, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h76, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he3, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h74, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h7c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h7e, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he9, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hea, 3'bzzz}: insn_immed_is_8bit = ~|(2'h3 & (2'b1 << immed_num));
    {8'heb, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hff, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hff, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h73, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h77, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h75, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h7d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h7f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h71, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h7b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h79, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h70, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h7a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h78, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h9f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc5, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc9, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc4, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hac, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'had, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he2, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he1, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he0, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h88, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h89, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc6, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc7, 3'h0}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hb0, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb1, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb2, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb3, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb4, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb5, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb6, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb7, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hb8, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hb9, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hba, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hbb, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hbc, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hbd, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hbe, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hbf, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h8e, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8e, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8e, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8e, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8e, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8e, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8e, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8e, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8c, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'ha0, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'ha1, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'ha2, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'ha3, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'ha4, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'ha5, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf6, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf7, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf6, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf7, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h90, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf6, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf7, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h08, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h09, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h0a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h0b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h0c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h0d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h1}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he6, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hee, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h6e, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h6f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'he7, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hef, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h58, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h59, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h5a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h5b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h5c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h5d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h5e, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h5f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h07, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h17, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h1f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h8f, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h61, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h9d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hff, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h06, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h0e, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h16, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h1e, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h50, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h51, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h52, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h53, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h54, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h55, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h56, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h57, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h68, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h6a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h60, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h9c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd0, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h2}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd0, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc3, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc2, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hcb, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hca, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hd0, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd0, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h9e, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd0, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd0, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h7}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h18, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h19, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h1a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h1b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h1c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h1d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h3}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h3}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hae, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'haf, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd6, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd0, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h4}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd0, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd1, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc0, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hc1, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd2, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd3, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf9, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hfd, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hfb, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'haa, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hab, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h28, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h29, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h2a, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h2b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h2c, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h2d, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h5}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h5}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h84, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h85, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'ha8, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'ha9, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hf6, 3'h0}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf6, 3'h1}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hf7, 3'h0}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'hf7, 3'h1}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h9b, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h86, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h87, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h91, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h92, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h93, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h94, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h95, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h96, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h97, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'hd7, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h30, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h31, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h32, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h33, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h34, 3'bzzz}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h35, 3'bzzz}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h80, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h81, 3'h6}: insn_immed_is_8bit = ~|(2'h1 & (2'b1 << immed_num));
    {8'h82, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    {8'h83, 3'h6}: insn_immed_is_8bit = ~|(2'h0 & (2'b1 << immed_num));
    default: insn_immed_is_8bit = 1'b0;
    endcase
endfunction
