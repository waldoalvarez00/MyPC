// Formal verification harness for FPU_RegisterStack
// Verifies stack pointer invariants, tag consistency, and overflow/underflow detection

`default_nettype none

module FPU_RegisterStack_formal (
    input logic clk
);
    // Reset signal
    logic reset;

    // Stack operations
    (* anyseq *) logic push;
    (* anyseq *) logic pop;
    (* anyseq *) logic inc_ptr;
    (* anyseq *) logic dec_ptr;
    (* anyseq *) logic free_reg;
    (* anyseq *) logic [2:0] free_index;
    (* anyseq *) logic init_stack;

    // Data interface
    (* anyseq *) logic [79:0] data_in;
    (* anyseq *) logic [2:0] write_reg;
    (* anyseq *) logic write_enable;
    (* anyseq *) logic [2:0] read_sel;

    // Outputs
    logic [79:0] st0, st1;
    logic [2:0] read_reg_out;
    logic [79:0] read_data;
    logic [2:0] stack_ptr;
    logic [15:0] tag_word;
    logic stack_overflow;
    logic stack_underflow;

    // Instantiate DUT
    FPU_RegisterStack dut (
        .clk(clk),
        .reset(reset),
        .push(push),
        .pop(pop),
        .inc_ptr(inc_ptr),
        .dec_ptr(dec_ptr),
        .free_reg(free_reg),
        .free_index(free_index),
        .init_stack(init_stack),
        .data_in(data_in),
        .write_reg(write_reg),
        .write_enable(write_enable),
        .st0(st0),
        .st1(st1),
        .read_reg(read_reg_out),
        .read_sel(read_sel),
        .read_data(read_data),
        .stack_ptr(stack_ptr),
        .tag_word(tag_word),
        .stack_overflow(stack_overflow),
        .stack_underflow(stack_underflow)
    );

    //=========================================================================
    // Reset sequence
    //=========================================================================

    logic seen_reset;

    initial begin
        reset = 1'b1;
        seen_reset = 1'b0;
    end

    always_ff @(posedge clk) begin
        if ($initstate) begin
            reset <= 1'b1;
            seen_reset <= 1'b0;
        end else begin
            reset <= 1'b0;
            if (reset)
                seen_reset <= 1'b1;
        end
    end

    //=========================================================================
    // Environment assumptions
    //=========================================================================

    // Only one stack operation at a time (realistic constraint)
    always_comb begin
        assume(!(push && pop));
        assume(!(push && inc_ptr));
        assume(!(push && dec_ptr));
        assume(!(pop && inc_ptr));
        assume(!(pop && dec_ptr));
        assume(!(inc_ptr && dec_ptr));
    end

    //=========================================================================
    // Shadow tracking for stack pointer
    //=========================================================================

    logic [2:0] shadow_sp;
    logic [2:0] expected_sp;

    always_ff @(posedge clk) begin
        if (reset) begin
            shadow_sp <= 3'd0;
        end else if (init_stack) begin
            shadow_sp <= 3'd0;
        end else begin
            expected_sp = shadow_sp;
            if (push)
                expected_sp = shadow_sp - 3'd1;
            else if (pop)
                expected_sp = shadow_sp + 3'd1;
            else if (inc_ptr)
                expected_sp = shadow_sp + 3'd1;
            else if (dec_ptr)
                expected_sp = shadow_sp - 3'd1;
            shadow_sp <= expected_sp;
        end
    end

    //=========================================================================
    // Formal Properties
    //=========================================================================

    always_ff @(posedge clk) begin
        if (seen_reset && !reset) begin

            //=================================================================
            // Property 1: Stack pointer always valid (implicitly 0-7 for 3 bits)
            //=================================================================
            // This is automatic for 3-bit value, but verify it tracks correctly
            assert(stack_ptr == shadow_sp);

            //=================================================================
            // Property 2: Init_stack resets stack pointer to 0
            //=================================================================
            if ($past(init_stack) && !$past(reset))
                assert(stack_ptr == 3'd0);

            //=================================================================
            // Property 3: Init_stack marks all registers as empty (tag = 11)
            //=================================================================
            if ($past(init_stack) && !$past(reset)) begin
                assert(tag_word[1:0] == 2'b11);    // ST(0)
                assert(tag_word[3:2] == 2'b11);    // ST(1)
                assert(tag_word[5:4] == 2'b11);    // ST(2)
                assert(tag_word[7:6] == 2'b11);    // ST(3)
                assert(tag_word[9:8] == 2'b11);    // ST(4)
                assert(tag_word[11:10] == 2'b11); // ST(5)
                assert(tag_word[13:12] == 2'b11); // ST(6)
                assert(tag_word[15:14] == 2'b11); // ST(7)
            end

            //=================================================================
            // Property 4: Push decrements stack pointer
            //=================================================================
            if ($past(push) && !$past(pop) && !$past(inc_ptr) && !$past(dec_ptr) &&
                !$past(init_stack) && !$past(reset))
                assert(stack_ptr == $past(stack_ptr) - 3'd1);

            //=================================================================
            // Property 5: Pop increments stack pointer
            //=================================================================
            if ($past(pop) && !$past(push) && !$past(inc_ptr) && !$past(dec_ptr) &&
                !$past(init_stack) && !$past(reset))
                assert(stack_ptr == $past(stack_ptr) + 3'd1);

            //=================================================================
            // Property 6: Inc_ptr increments stack pointer (FINCSTP)
            //=================================================================
            if ($past(inc_ptr) && !$past(push) && !$past(pop) && !$past(dec_ptr) &&
                !$past(init_stack) && !$past(reset))
                assert(stack_ptr == $past(stack_ptr) + 3'd1);

            //=================================================================
            // Property 7: Dec_ptr decrements stack pointer (FDECSTP)
            //=================================================================
            if ($past(dec_ptr) && !$past(push) && !$past(pop) && !$past(inc_ptr) &&
                !$past(init_stack) && !$past(reset))
                assert(stack_ptr == $past(stack_ptr) - 3'd1);

            //=================================================================
            // Property 8: Overflow flag only asserted when pushing to non-empty
            //=================================================================
            // If overflow is asserted, push must have occurred
            if (stack_overflow)
                assert($past(push));

            //=================================================================
            // Property 9: Underflow flag only asserted when popping from empty
            //=================================================================
            // If underflow is asserted, pop must have occurred
            if (stack_underflow)
                assert($past(pop));

            //=================================================================
            // Property 10: Free_reg marks register as empty
            //=================================================================
            // After free_reg, the corresponding tag should be empty (11)
            // Note: This is complex due to physical_reg mapping, simplified check

            //=================================================================
            // Property 11: No spurious overflow/underflow on reset
            //=================================================================
            if ($past(reset)) begin
                assert(!stack_overflow);
                assert(!stack_underflow);
            end

            //=================================================================
            // Property 12: Tag word correctly reflects empty on init
            //=================================================================
            // After reset, all tags should be empty
            if ($fell(reset)) begin
                assert(tag_word == 16'hFFFF);  // All 11s
            end

        end
    end

    //=========================================================================
    // Cover Properties - Verify reachability
    //=========================================================================

    always_ff @(posedge clk) begin
        if (seen_reset && !reset) begin
            // Cover: Stack overflow occurs
            cover(stack_overflow);

            // Cover: Stack underflow occurs
            cover(stack_underflow);

            // Cover: Push operation
            cover(push && !pop);

            // Cover: Pop operation
            cover(pop && !push);

            // Cover: Free register
            cover(free_reg);

            // Cover: Init stack
            cover(init_stack);

            // Cover: Write to register
            cover(write_enable);

            // Cover: Stack pointer wraps around (7 -> 0)
            cover(stack_ptr == 3'd0 && $past(stack_ptr) == 3'd7);

            // Cover: Stack pointer wraps around (0 -> 7)
            cover(stack_ptr == 3'd7 && $past(stack_ptr) == 3'd0);

            // Cover: Various stack pointer values
            cover(stack_ptr == 3'd0);
            cover(stack_ptr == 3'd4);
            cover(stack_ptr == 3'd7);
        end
    end

endmodule
