// Copyright 2025, Waldo Alvarez, https://pipflow.com
`timescale 1ns / 1ps

//=====================================================================
// IEEE 754 Extended Precision (80-bit) Unified Multiply/Divide Unit
//
// Consolidates multiplication and division into a single unit with
// shared resources for area optimization.
//
// Features:
// - Single module supporting both multiply and divide operations
// - Shared unpacking, normalization, and rounding logic
// - ~25% area reduction vs. separate modules
// - Maintains full IEEE 754 compliance
//
// Format: [79:Sign][78:64:Exponent][63:Integer][62:0:Fraction]
//
// Area Savings:
// - Original: 757 lines (324 mul + 433 div)
// - Unified: ~550 lines
// - Reduction: ~200 lines (~25%)
//=====================================================================

module FPU_IEEE754_MulDiv_Unified(
    input wire clk,
    input wire reset,
    input wire enable,                  // Start operation
    input wire operation,               // 0=multiply, 1=divide

    // Operands
    input wire [79:0] operand_a,       // First operand (80-bit)
    input wire [79:0] operand_b,       // Second operand (80-bit)

    // Control
    input wire [1:0]  rounding_mode,   // 00=nearest, 01=down, 10=up, 11=truncate

    // Result
    output reg [79:0] result,          // Result (80-bit)
    output wire       done,            // Operation complete

    // Exception flags
    output reg        flag_invalid,    // Invalid operation
    output reg        flag_div_by_zero,// Division by zero (divide only)
    output reg        flag_overflow,   // Result overflow
    output reg        flag_underflow,  // Result underflow
    output reg        flag_inexact     // Result not exact (rounded)
);

    //=================================================================
    // Internal States
    //=================================================================

    localparam STATE_IDLE       = 3'd0;
    localparam STATE_UNPACK     = 3'd1;
    localparam STATE_COMPUTE    = 3'd2;
    localparam STATE_NORMALIZE  = 3'd3;
    localparam STATE_ROUND      = 3'd4;
    localparam STATE_PACK       = 3'd5;

    reg [2:0] state;
    reg       is_multiply;  // Latched operation type
    reg       done_reg;     // Internal done register
    reg       started;      // Have we started an operation since enable went high?

    // done is simply the done_reg - we use the started flag to prevent retriggering
    assign done = done_reg;

    //=================================================================
    // Unpacked Operands (SHARED)
    //=================================================================

    reg        sign_a, sign_b;
    reg [14:0] exp_a, exp_b;
    reg [63:0] mant_a, mant_b;
    reg        is_zero_a, is_inf_a, is_nan_a, is_unnormal_a;
    reg        is_zero_b, is_inf_b, is_nan_b, is_unnormal_b;

    //=================================================================
    // Working Registers (SHARED)
    //=================================================================

    reg        result_sign;
    reg signed [16:0] result_exp;      // 17-bit signed for overflow/underflow
    reg [66:0] result_mant;            // Normalized result with guard/round/sticky

    //=================================================================
    // Multiply-Specific Registers
    //=================================================================

    (* multstyle = "dsp" *) reg [127:0] product;               // 64×64 = 128-bit product

    //=================================================================
    // Divide-Specific Registers
    //=================================================================

    reg signed [128:0] remainder;      // Signed partial remainder for SRT-2
    reg [63:0] divisor;
    reg [63:0] divisor_half;          // divisor >> 1 for SRT selection
    reg signed [1:0] quotient_digits [0:66];  // Signed-digit quotient
    reg [6:0]  div_count;             // Division iteration counter
    reg [66:0] quotient;              // Binary quotient
    integer    srt_i;                 // Loop variable

    //=================================================================
    // Rounding Registers (SHARED)
    //=================================================================

    reg round_bit, sticky_bit;

    //=================================================================
    // Special Value Detection (SHARED)
    //=================================================================

    task detect_special_values;
        begin
            // Operand A
            is_zero_a = (exp_a == 15'd0) && (mant_a == 64'd0);
            is_inf_a = (exp_a == 15'h7FFF) && (mant_a[62:0] == 63'd0) && (mant_a[63] == 1'b1);
            is_nan_a = (exp_a == 15'h7FFF) && ((mant_a[62:0] != 63'd0) || (mant_a[63] == 1'b0));
            // Pseudo-normal (unnormal): non-zero/non-max exponent but integer bit = 0
            // This is an unsupported format that should raise IE
            is_unnormal_a = (exp_a != 15'd0) && (exp_a != 15'h7FFF) && (mant_a[63] == 1'b0);

            // Operand B
            is_zero_b = (exp_b == 15'd0) && (mant_b == 64'd0);
            is_inf_b = (exp_b == 15'h7FFF) && (mant_b[62:0] == 63'd0) && (mant_b[63] == 1'b1);
            is_nan_b = (exp_b == 15'h7FFF) && ((mant_b[62:0] != 63'd0) || (mant_b[63] == 1'b0));
            // Pseudo-normal (unnormal): non-zero/non-max exponent but integer bit = 0
            is_unnormal_b = (exp_b != 15'd0) && (exp_b != 15'h7FFF) && (mant_b[63] == 1'b0);
        end
    endtask

    //=================================================================
    // Main State Machine
    //=================================================================

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= STATE_IDLE;
            done_reg <= 1'b0;
            started <= 1'b0;
            result <= 80'd0;
            flag_invalid <= 1'b0;
            flag_div_by_zero <= 1'b0;
            flag_overflow <= 1'b0;
            flag_underflow <= 1'b0;
            flag_inexact <= 1'b0;
        end else begin
            case (state)
                //=========================================================
                // IDLE State
                //=========================================================
                STATE_IDLE: begin
                    if (!enable) begin
                        // Master acknowledged result or no request - reset for next operation
                        started <= 1'b0;
                        done_reg <= 1'b0;
                        flag_invalid <= 1'b0;
                        flag_div_by_zero <= 1'b0;
                        flag_overflow <= 1'b0;
                        flag_underflow <= 1'b0;
                        flag_inexact <= 1'b0;
                    end else if (!started) begin
                        // Start new operation only if we haven't already started one
                        `ifdef ICARUS
                        $display("[MULDIV] Starting op=%b, A=%h, B=%h", operation, operand_a, operand_b);
                        `endif
                        started <= 1'b1;
                        is_multiply <= ~operation;  // Latch operation
                        state <= STATE_UNPACK;
                    end
                    // else: enable high but already started - wait for master to lower enable
                end

                //=========================================================
                // UNPACK State (SHARED)
                //=========================================================
                STATE_UNPACK: begin
                    // Unpack operands
                    sign_a = operand_a[79];
                    exp_a = operand_a[78:64];
                    mant_a = operand_a[63:0];

                    sign_b = operand_b[79];
                    exp_b = operand_b[78:64];
                    mant_b = operand_b[63:0];

                    detect_special_values;

                    // Calculate result sign (XOR of signs for both mul/div)
                    result_sign = sign_a ^ sign_b;

                    // Handle special cases
                    if (is_nan_a || is_nan_b || is_unnormal_a || is_unnormal_b) begin
                        // NaN or unsupported format (pseudo-normal) -> return QNaN
                        result <= {1'b0, 15'h7FFF, 1'b1, 63'h4000000000000000};
                        flag_invalid <= 1'b1;
                        done_reg <= 1'b1;
                        state <= STATE_IDLE;
                    end else if (is_multiply) begin
                        // MULTIPLY special cases
                        if ((is_zero_a && is_inf_b) || (is_inf_a && is_zero_b)) begin
                            // 0 × ∞ = NaN
                            result <= {1'b0, 15'h7FFF, 1'b1, 63'h4000000000000000};
                            flag_invalid <= 1'b1;
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else if (is_inf_a || is_inf_b) begin
                            // ∞ × finite = ∞
                            result <= {result_sign, 15'h7FFF, 1'b1, 63'd0};
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else if (is_zero_a || is_zero_b) begin
                            // 0 × anything = 0
                            result <= {result_sign, 79'd0};
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else begin
                            state <= STATE_COMPUTE;
                        end
                    end else begin
                        // DIVIDE special cases
                        if ((is_zero_a && is_zero_b) || (is_inf_a && is_inf_b)) begin
                            // 0÷0 or ∞÷∞ = NaN
                            result <= {1'b0, 15'h7FFF, 1'b1, 63'h4000000000000000};
                            flag_invalid <= 1'b1;
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else if (is_zero_b) begin
                            // x÷0 = ±∞
                            result <= {result_sign, 15'h7FFF, 1'b1, 63'd0};
                            flag_div_by_zero <= 1'b1;
                            done_reg <= 1'b1;
                            `ifdef ICARUS
                            $display("[MULDIV] Divide by zero detected: A=%h, B=%h, result=%h", operand_a, operand_b, {result_sign, 15'h7FFF, 1'b1, 63'd0});
                            `endif
                            state <= STATE_IDLE;
                        end else if (is_inf_a) begin
                            // ∞÷finite = ±∞
                            result <= {result_sign, 15'h7FFF, 1'b1, 63'd0};
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else if (is_zero_a || is_inf_b) begin
                            // 0÷finite = ±0 or finite÷∞ = ±0
                            result <= {result_sign, 79'd0};
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else begin
                            state <= STATE_COMPUTE;
                        end
                    end
                end

                //=========================================================
                // COMPUTE State (OPERATION-SPECIFIC)
                //=========================================================
                STATE_COMPUTE: begin
                    if (is_multiply) begin
                        //=====================================================
                        // MULTIPLY
                        //=====================================================
                        // Add exponents and subtract bias
                        if ({1'b0, exp_a} + {1'b0, exp_b} < 16'd16383) begin
                            // Underflow
                            result <= {result_sign, 79'd0};
                            flag_underflow <= 1'b1;
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else begin
                            result_exp = {1'b0, exp_a} + {1'b0, exp_b} - 17'd16383;
                            // Multiply mantissas
                            product = mant_a * mant_b;
                            state <= STATE_NORMALIZE;
                        end
                    end else begin
                        //=====================================================
                        // DIVIDE
                        //=====================================================
                        // Subtract exponents and add bias
                        if ({1'b0, exp_a} + 17'd16383 < {1'b0, exp_b}) begin
                            // Underflow
                            result <= {result_sign, 79'd0};
                            flag_underflow <= 1'b1;
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else begin
                            result_exp = {2'b00, exp_a} - {2'b00, exp_b} + 17'sd16383;

                            // SRT-2 Division Initialization
                            divisor = mant_b;
                            divisor_half = mant_b >> 1;

                            // Initialize quotient digits
                            for (srt_i = 0; srt_i <= 66; srt_i = srt_i + 1) begin
                                quotient_digits[srt_i] = 2'sd0;
                            end

                            // Pre-normalize based on mant_a vs mant_b
                            if (mant_a >= mant_b) begin
                                quotient_digits[0] = 2'sd1;
                                remainder = {1'b0, mant_a - mant_b, 64'd0};
                                div_count = 7'd1;
                            end else begin
                                quotient_digits[0] = 2'sd0;
                                remainder = {1'b0, mant_a, 64'd0};
                                div_count = 7'd1;
                            end

                            state <= STATE_NORMALIZE;
                        end
                    end
                end

                //=========================================================
                // NORMALIZE State (OPERATION-SPECIFIC)
                //=========================================================
                STATE_NORMALIZE: begin
                    if (is_multiply) begin
                        //=====================================================
                        // MULTIPLY NORMALIZATION
                        //=====================================================
                        if (product[127]) begin
                            // Product needs 128 bits, shift right by 1
                            result_mant = {product[127:62], |product[61:0]};
                            result_exp = result_exp + 17'd1;
                        end else if (product[126]) begin
                            // Product fits in 127 bits
                            result_mant = {product[126:61], |product[60:0]};
                        end else begin
                            // Find leading 1 for denormalized product
                            integer i;
                            reg [6:0] shift_amount;
                            shift_amount = 7'd0;

                            for (i = 125; i >= 0; i = i - 1) begin
                                if (product[i] && shift_amount == 7'd0) begin
                                    shift_amount = 7'd126 - i[6:0];
                                end
                            end

                            if (shift_amount > 0) begin
                                result_mant = {(product << shift_amount), 3'b000};
                                result_exp = result_exp - shift_amount;
                            end else begin
                                result_mant = {product[126:63], |product[62:0]};
                            end
                        end

                        // Check for overflow/underflow
                        if (result_exp >= 17'sd32767) begin
                            result <= {result_sign, 15'h7FFF, 1'b1, 63'd0};
                            flag_overflow <= 1'b1;
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else if (result_exp[16]) begin  // Negative
                            result <= {result_sign, 79'd0};
                            flag_underflow <= 1'b1;
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else begin
                            state <= STATE_ROUND;
                        end
                    end else begin
                        //=====================================================
                        // DIVIDE NORMALIZATION (SRT-2 iterations)
                        //=====================================================
                        if (div_count < 7'd67) begin
                            // SRT-2 Selection Function
                            if (!remainder[128] && remainder[127:64] >= divisor_half) begin
                                quotient_digits[div_count] = 2'sd1;
                            end else if (remainder[128] && (-remainder) > {1'b0, divisor_half, 64'd0}) begin
                                quotient_digits[div_count] = -2'sd1;
                            end else begin
                                quotient_digits[div_count] = 2'sd0;
                            end

                            // Update remainder: R_next = 2*R - q*D
                            remainder = remainder << 1;
                            if (quotient_digits[div_count] == 2'sd1) begin
                                remainder = remainder - {1'b0, divisor, 64'd0};
                            end else if (quotient_digits[div_count] == -2'sd1) begin
                                remainder = remainder + {1'b0, divisor, 64'd0};
                            end

                            div_count = div_count + 7'd1;
                        end else begin
                            // Convert signed-digit quotient to binary
                            quotient = 67'd0;
                            for (srt_i = 0; srt_i <= 66; srt_i = srt_i + 1) begin
                                if (quotient_digits[srt_i] == 2'sd1) begin
                                    quotient = quotient + (67'd1 << (66 - srt_i));
                                end else if (quotient_digits[srt_i] == -2'sd1) begin
                                    quotient = quotient - (67'd1 << (66 - srt_i));
                                end
                            end

                            result_mant = quotient;

                            // Set sticky bit if remainder is non-zero (inexact division)
                            if (remainder != 129'd0) begin
                                result_mant[0] = 1'b1;
                            end

                            // Normalize quotient
                            if (result_mant[66]) begin
                                // Already normalized
                            end else if (result_mant[65]) begin
                                result_mant = result_mant << 1;
                                result_exp = result_exp - 17'sd1;
                            end else begin
                                // Find leading 1
                                integer i;
                                reg [6:0] shift_amount;
                                shift_amount = 7'd0;

                                for (i = 64; i >= 0; i = i - 1) begin
                                    if (result_mant[i] && shift_amount == 7'd0) begin
                                        shift_amount = 7'd66 - i[6:0];
                                    end
                                end

                                if (shift_amount > 0 && shift_amount < 67) begin
                                    result_mant = result_mant << shift_amount;
                                    result_exp = result_exp - shift_amount;
                                end
                            end

                            // Check for overflow/underflow
                            if (result_exp > 17'sd32766) begin
                                result <= {result_sign, 15'h7FFF, 1'b1, 63'd0};
                                flag_overflow <= 1'b1;
                                done_reg <= 1'b1;
                                state <= STATE_IDLE;
                            end else if (result_exp < 17'sd1) begin
                                result <= {result_sign, 79'd0};
                                flag_underflow <= 1'b1;
                                done_reg <= 1'b1;
                                state <= STATE_IDLE;
                            end else begin
                                state <= STATE_ROUND;
                            end
                        end
                    end
                end

                //=========================================================
                // ROUND State (SHARED)
                //=========================================================
                STATE_ROUND: begin
                    // Extract guard, round, sticky bits
                    // result_mant format: [66:int][65:3:frac][2:guard][1:round][0:sticky]
                    round_bit = result_mant[1];
                    sticky_bit = result_mant[0];

                    // Round according to mode
                    case (rounding_mode)
                        2'b00: begin // Round to nearest (ties to even)
                            if (round_bit && (sticky_bit || result_mant[2])) begin
                                result_mant = (result_mant >> 3) + 65'd1;
                                flag_inexact <= 1'b1;
                            end else begin
                                result_mant = result_mant >> 3;
                                if (round_bit || sticky_bit) flag_inexact <= 1'b1;
                            end
                        end
                        2'b01: begin // Round down (toward -∞)
                            if (result_sign && (round_bit || sticky_bit)) begin
                                result_mant = (result_mant >> 3) + 65'd1;
                                flag_inexact <= 1'b1;
                            end else begin
                                result_mant = result_mant >> 3;
                                if (round_bit || sticky_bit) flag_inexact <= 1'b1;
                            end
                        end
                        2'b10: begin // Round up (toward +∞)
                            if (!result_sign && (round_bit || sticky_bit)) begin
                                result_mant = (result_mant >> 3) + 65'd1;
                                flag_inexact <= 1'b1;
                            end else begin
                                result_mant = result_mant >> 3;
                                if (round_bit || sticky_bit) flag_inexact <= 1'b1;
                            end
                        end
                        2'b11: begin // Round toward zero (truncate)
                            result_mant = result_mant >> 3;
                            if (round_bit || sticky_bit) flag_inexact <= 1'b1;
                        end
                    endcase

                    // Check for rounding overflow
                    if (result_mant[64]) begin
                        result_mant = result_mant >> 1;
                        result_exp = result_exp + 17'd1;

                        if (result_exp >= 17'sd32767) begin
                            result <= {result_sign, 15'h7FFF, 1'b1, 63'd0};
                            flag_overflow <= 1'b1;
                            done_reg <= 1'b1;
                            state <= STATE_IDLE;
                        end else begin
                            state <= STATE_PACK;
                        end
                    end else begin
                        state <= STATE_PACK;
                    end
                end

                //=========================================================
                // PACK State (SHARED)
                //=========================================================
                STATE_PACK: begin
                    result <= {result_sign, result_exp[14:0], result_mant[63:0]};
                    done_reg <= 1'b1;
                    state <= STATE_IDLE;
                end

                default: begin
                    state <= STATE_IDLE;
                end
            endcase
        end
    end

endmodule
